// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_clk,         // alt_vip_cl_cvo_hdmi_clocked_video.vid_clk
		output wire [31:0] alt_vip_cl_cvo_hdmi_clocked_video_vid_data,        //                                  .vid_data
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_underflow,       //                                  .underflow
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_mode_change, //                                  .vid_mode_change
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_std,         //                                  .vid_std
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_datavalid,   //                                  .vid_datavalid
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_v_sync,      //                                  .vid_v_sync
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_h_sync,      //                                  .vid_h_sync
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_f,           //                                  .vid_f
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_h,           //                                  .vid_h
		output wire        alt_vip_cl_cvo_hdmi_clocked_video_vid_v,           //                                  .vid_v
		inout  wire [7:0]  arduino_gpio_export,                               //                      arduino_gpio.export
		input  wire [1:0]  button_pio_export,                                 //                        button_pio.export
		input  wire        clk_clk,                                           //                               clk.clk
		output wire        clk_hdmi_clk,                                      //                          clk_hdmi.clk
		output wire [1:0]  ctrl_reg_export,                                   //                          ctrl_reg.export
		input  wire [3:0]  dipsw_pio_export,                                  //                         dipsw_pio.export
		inout  wire [17:0] gpio_0_a_export,                                   //                          gpio_0_a.export
		inout  wire [17:0] gpio_0_b_export,                                   //                          gpio_0_b.export
		inout  wire [17:0] gpio_1_a_export,                                   //                          gpio_1_a.export
		inout  wire [17:0] gpio_1_b_export,                                   //                          gpio_1_b.export
		input  wire        hps_0_f2h_cold_reset_req_reset_n,                  //          hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,                 //         hps_0_f2h_debug_reset_req.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,              //           hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,                  //          hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,                           //                   hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,             //                      hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,               //                                  .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,               //                                  .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,               //                                  .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,               //                                  .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,               //                                  .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,               //                                  .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,                //                                  .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,             //                                  .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,             //                                  .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,             //                                  .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,               //                                  .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,               //                                  .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,               //                                  .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,                 //                                  .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,                  //                                  .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,                  //                                  .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,                 //                                  .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,                  //                                  .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,                  //                                  .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,                  //                                  .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,                  //                                  .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,                  //                                  .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,                  //                                  .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,                  //                                  .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,                  //                                  .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,                  //                                  .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,                  //                                  .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,                 //                                  .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,                 //                                  .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,                 //                                  .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,                 //                                  .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,                //                                  .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,               //                                  .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,               //                                  .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,                //                                  .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,                 //                                  .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,                 //                                  .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,                 //                                  .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,                 //                                  .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,                 //                                  .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,                 //                                  .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,              //                                  .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,              //                                  .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,              //                                  .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,              //                                  .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,              //                                  .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,              //                                  .hps_io_gpio_inst_GPIO61
		output wire        hps_0_i2c2_out_data,                               //                        hps_0_i2c2.out_data
		input  wire        hps_0_i2c2_sda,                                    //                                  .sda
		output wire        hps_0_i2c2_clk_clk,                                //                    hps_0_i2c2_clk.clk
		input  wire        hps_0_i2c2_scl_in_clk,                             //                 hps_0_i2c2_scl_in.clk
		output wire        hps_0_i2c3_out_data,                               //                        hps_0_i2c3.out_data
		input  wire        hps_0_i2c3_sda,                                    //                                  .sda
		output wire        hps_0_i2c3_clk_clk,                                //                    hps_0_i2c3_clk.clk
		input  wire        hps_0_i2c3_scl_in_clk,                             //                 hps_0_i2c3_scl_in.clk
		output wire        hps_0_spim0_txd,                                   //                       hps_0_spim0.txd
		input  wire        hps_0_spim0_rxd,                                   //                                  .rxd
		input  wire        hps_0_spim0_ss_in_n,                               //                                  .ss_in_n
		output wire        hps_0_spim0_ssi_oe_n,                              //                                  .ssi_oe_n
		output wire        hps_0_spim0_ss_0_n,                                //                                  .ss_0_n
		output wire        hps_0_spim0_ss_1_n,                                //                                  .ss_1_n
		output wire        hps_0_spim0_ss_2_n,                                //                                  .ss_2_n
		output wire        hps_0_spim0_ss_3_n,                                //                                  .ss_3_n
		output wire        hps_0_spim0_sclk_out_clk,                          //              hps_0_spim0_sclk_out.clk
		input  wire        hps_0_uart1_cts,                                   //                       hps_0_uart1.cts
		input  wire        hps_0_uart1_dsr,                                   //                                  .dsr
		input  wire        hps_0_uart1_dcd,                                   //                                  .dcd
		input  wire        hps_0_uart1_ri,                                    //                                  .ri
		output wire        hps_0_uart1_dtr,                                   //                                  .dtr
		output wire        hps_0_uart1_rts,                                   //                                  .rts
		output wire        hps_0_uart1_out1_n,                                //                                  .out1_n
		output wire        hps_0_uart1_out2_n,                                //                                  .out2_n
		input  wire        hps_0_uart1_rxd,                                   //                                  .rxd
		output wire        hps_0_uart1_txd,                                   //                                  .txd
		output wire [7:0]  led_pio_export,                                    //                           led_pio.export
		output wire [14:0] memory_mem_a,                                      //                            memory.mem_a
		output wire [2:0]  memory_mem_ba,                                     //                                  .mem_ba
		output wire        memory_mem_ck,                                     //                                  .mem_ck
		output wire        memory_mem_ck_n,                                   //                                  .mem_ck_n
		output wire        memory_mem_cke,                                    //                                  .mem_cke
		output wire        memory_mem_cs_n,                                   //                                  .mem_cs_n
		output wire        memory_mem_ras_n,                                  //                                  .mem_ras_n
		output wire        memory_mem_cas_n,                                  //                                  .mem_cas_n
		output wire        memory_mem_we_n,                                   //                                  .mem_we_n
		output wire        memory_mem_reset_n,                                //                                  .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                     //                                  .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                    //                                  .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                  //                                  .mem_dqs_n
		output wire        memory_mem_odt,                                    //                                  .mem_odt
		output wire [3:0]  memory_mem_dm,                                     //                                  .mem_dm
		input  wire        memory_oct_rzqin,                                  //                                  .oct_rzqin
		input  wire [31:0] random_reg_export,                                 //                        random_reg.export
		output wire [31:0] reset_val_export                                   //                         reset_val.export
	);

	wire          alt_vip_cl_vfb_hdmi_dout_valid;                                      // alt_vip_cl_vfb_hdmi:dout_valid -> alt_vip_cl_cvo_hdmi:din_valid
	wire   [31:0] alt_vip_cl_vfb_hdmi_dout_data;                                       // alt_vip_cl_vfb_hdmi:dout_data -> alt_vip_cl_cvo_hdmi:din_data
	wire          alt_vip_cl_vfb_hdmi_dout_ready;                                      // alt_vip_cl_cvo_hdmi:din_ready -> alt_vip_cl_vfb_hdmi:dout_ready
	wire          alt_vip_cl_vfb_hdmi_dout_startofpacket;                              // alt_vip_cl_vfb_hdmi:dout_startofpacket -> alt_vip_cl_cvo_hdmi:din_startofpacket
	wire          alt_vip_cl_vfb_hdmi_dout_endofpacket;                                // alt_vip_cl_vfb_hdmi:dout_endofpacket -> alt_vip_cl_cvo_hdmi:din_endofpacket
	wire          hps_0_h2f_user0_clock_clk;                                           // hps_0:h2f_user0_clk -> [alt_vip_cl_vfb_hdmi:mem_clock, hps_0:f2h_axi_clk, hps_0:f2h_sdram0_clk, mm_interconnect_5:hps_0_h2f_user0_clock_clk, rst_controller:clk, rst_controller_006:clk]
	wire          hps_0_h2f_user1_clock_clk;                                           // hps_0:h2f_user1_clk -> rst_controller_004:clk
	wire          pll_stream_outclk0_clk;                                              // pll_stream:outclk_0 -> custom_reset_synchronizer:clk_in
	wire          pll_reset_pio_external_connection_export;                            // pll_reset_pio:out_port -> pll_stream:rst
	wire          cvo_reset_pio_external_connection_export;                            // cvo_reset_pio:out_port -> rst_controller_003:reset_in1
	wire          pll_stream_locked_export;                                            // pll_stream:locked -> locked_pio:in_port
	wire   [63:0] pll_stream_reconfig_from_pll_reconfig_from_pll;                      // pll_stream:reconfig_from_pll -> pll_stream_reconfig:reconfig_from_pll
	wire   [63:0] pll_stream_reconfig_reconfig_to_pll_reconfig_to_pll;                 // pll_stream_reconfig:reconfig_to_pll -> pll_stream:reconfig_to_pll
	wire          custom_reset_synchronizer_reset_out_reset;                           // custom_reset_synchronizer:reset_out -> [alt_vip_cl_cvo_hdmi:main_reset_reset, alt_vip_cl_vfb_hdmi:main_reset, hdmi_mm_bridge:reset, mm_interconnect_2:hdmi_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_3:hdmi_mm_bridge_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0]
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                        // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                          // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                          // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                         // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                            // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                         // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                          // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                            // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                        // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                         // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                         // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                         // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                         // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                          // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                        // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                        // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                           // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                         // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                         // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                         // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                          // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                        // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                          // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                        // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                        // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                         // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                         // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                          // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                          // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                          // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                           // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                            // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                         // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                         // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                        // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                         // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [31:0] mm_interconnect_0_custom_ip_bridge_s0_readdata;                      // custom_ip_bridge:s0_readdata -> mm_interconnect_0:custom_ip_bridge_s0_readdata
	wire          mm_interconnect_0_custom_ip_bridge_s0_waitrequest;                   // custom_ip_bridge:s0_waitrequest -> mm_interconnect_0:custom_ip_bridge_s0_waitrequest
	wire          mm_interconnect_0_custom_ip_bridge_s0_debugaccess;                   // mm_interconnect_0:custom_ip_bridge_s0_debugaccess -> custom_ip_bridge:s0_debugaccess
	wire    [5:0] mm_interconnect_0_custom_ip_bridge_s0_address;                       // mm_interconnect_0:custom_ip_bridge_s0_address -> custom_ip_bridge:s0_address
	wire          mm_interconnect_0_custom_ip_bridge_s0_read;                          // mm_interconnect_0:custom_ip_bridge_s0_read -> custom_ip_bridge:s0_read
	wire    [3:0] mm_interconnect_0_custom_ip_bridge_s0_byteenable;                    // mm_interconnect_0:custom_ip_bridge_s0_byteenable -> custom_ip_bridge:s0_byteenable
	wire          mm_interconnect_0_custom_ip_bridge_s0_readdatavalid;                 // custom_ip_bridge:s0_readdatavalid -> mm_interconnect_0:custom_ip_bridge_s0_readdatavalid
	wire          mm_interconnect_0_custom_ip_bridge_s0_write;                         // mm_interconnect_0:custom_ip_bridge_s0_write -> custom_ip_bridge:s0_write
	wire   [31:0] mm_interconnect_0_custom_ip_bridge_s0_writedata;                     // mm_interconnect_0:custom_ip_bridge_s0_writedata -> custom_ip_bridge:s0_writedata
	wire    [0:0] mm_interconnect_0_custom_ip_bridge_s0_burstcount;                    // mm_interconnect_0:custom_ip_bridge_s0_burstcount -> custom_ip_bridge:s0_burstcount
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;                    // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                      // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                       // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire    [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                    // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;                         // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                     // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;                         // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                     // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                       // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                       // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                      // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                       // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                         // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                     // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                      // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                      // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                      // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                      // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                       // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                     // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                     // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                        // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                      // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                      // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                      // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                     // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                     // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                      // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                      // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                       // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                        // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                      // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                     // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                      // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] mm_interconnect_1_lw_mm_bridge_s0_readdata;                          // lw_mm_bridge:s0_readdata -> mm_interconnect_1:lw_mm_bridge_s0_readdata
	wire          mm_interconnect_1_lw_mm_bridge_s0_waitrequest;                       // lw_mm_bridge:s0_waitrequest -> mm_interconnect_1:lw_mm_bridge_s0_waitrequest
	wire          mm_interconnect_1_lw_mm_bridge_s0_debugaccess;                       // mm_interconnect_1:lw_mm_bridge_s0_debugaccess -> lw_mm_bridge:s0_debugaccess
	wire   [16:0] mm_interconnect_1_lw_mm_bridge_s0_address;                           // mm_interconnect_1:lw_mm_bridge_s0_address -> lw_mm_bridge:s0_address
	wire          mm_interconnect_1_lw_mm_bridge_s0_read;                              // mm_interconnect_1:lw_mm_bridge_s0_read -> lw_mm_bridge:s0_read
	wire    [3:0] mm_interconnect_1_lw_mm_bridge_s0_byteenable;                        // mm_interconnect_1:lw_mm_bridge_s0_byteenable -> lw_mm_bridge:s0_byteenable
	wire          mm_interconnect_1_lw_mm_bridge_s0_readdatavalid;                     // lw_mm_bridge:s0_readdatavalid -> mm_interconnect_1:lw_mm_bridge_s0_readdatavalid
	wire          mm_interconnect_1_lw_mm_bridge_s0_write;                             // mm_interconnect_1:lw_mm_bridge_s0_write -> lw_mm_bridge:s0_write
	wire   [31:0] mm_interconnect_1_lw_mm_bridge_s0_writedata;                         // mm_interconnect_1:lw_mm_bridge_s0_writedata -> lw_mm_bridge:s0_writedata
	wire    [0:0] mm_interconnect_1_lw_mm_bridge_s0_burstcount;                        // mm_interconnect_1:lw_mm_bridge_s0_burstcount -> lw_mm_bridge:s0_burstcount
	wire          lw_mm_bridge_m0_waitrequest;                                         // mm_interconnect_2:lw_mm_bridge_m0_waitrequest -> lw_mm_bridge:m0_waitrequest
	wire   [31:0] lw_mm_bridge_m0_readdata;                                            // mm_interconnect_2:lw_mm_bridge_m0_readdata -> lw_mm_bridge:m0_readdata
	wire          lw_mm_bridge_m0_debugaccess;                                         // lw_mm_bridge:m0_debugaccess -> mm_interconnect_2:lw_mm_bridge_m0_debugaccess
	wire   [16:0] lw_mm_bridge_m0_address;                                             // lw_mm_bridge:m0_address -> mm_interconnect_2:lw_mm_bridge_m0_address
	wire          lw_mm_bridge_m0_read;                                                // lw_mm_bridge:m0_read -> mm_interconnect_2:lw_mm_bridge_m0_read
	wire    [3:0] lw_mm_bridge_m0_byteenable;                                          // lw_mm_bridge:m0_byteenable -> mm_interconnect_2:lw_mm_bridge_m0_byteenable
	wire          lw_mm_bridge_m0_readdatavalid;                                       // mm_interconnect_2:lw_mm_bridge_m0_readdatavalid -> lw_mm_bridge:m0_readdatavalid
	wire   [31:0] lw_mm_bridge_m0_writedata;                                           // lw_mm_bridge:m0_writedata -> mm_interconnect_2:lw_mm_bridge_m0_writedata
	wire          lw_mm_bridge_m0_write;                                               // lw_mm_bridge:m0_write -> mm_interconnect_2:lw_mm_bridge_m0_write
	wire    [0:0] lw_mm_bridge_m0_burstcount;                                          // lw_mm_bridge:m0_burstcount -> mm_interconnect_2:lw_mm_bridge_m0_burstcount
	wire          mm_interconnect_2_jtag_uart_avalon_jtag_slave_chipselect;            // mm_interconnect_2:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_2_jtag_uart_avalon_jtag_slave_readdata;              // jtag_uart:av_readdata -> mm_interconnect_2:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_2_jtag_uart_avalon_jtag_slave_waitrequest;           // jtag_uart:av_waitrequest -> mm_interconnect_2:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_2_jtag_uart_avalon_jtag_slave_address;               // mm_interconnect_2:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_2_jtag_uart_avalon_jtag_slave_read;                  // mm_interconnect_2:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_2_jtag_uart_avalon_jtag_slave_write;                 // mm_interconnect_2:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_2_jtag_uart_avalon_jtag_slave_writedata;             // mm_interconnect_2:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [31:0] mm_interconnect_2_sysid_qsys_control_slave_readdata;                 // sysid_qsys:readdata -> mm_interconnect_2:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_2_sysid_qsys_control_slave_address;                  // mm_interconnect_2:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_readdata;    // pll_stream_reconfig:mgmt_readdata -> mm_interconnect_2:pll_stream_reconfig_mgmt_avalon_slave_readdata
	wire          mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_waitrequest; // pll_stream_reconfig:mgmt_waitrequest -> mm_interconnect_2:pll_stream_reconfig_mgmt_avalon_slave_waitrequest
	wire    [5:0] mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_address;     // mm_interconnect_2:pll_stream_reconfig_mgmt_avalon_slave_address -> pll_stream_reconfig:mgmt_address
	wire          mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_read;        // mm_interconnect_2:pll_stream_reconfig_mgmt_avalon_slave_read -> pll_stream_reconfig:mgmt_read
	wire    [3:0] mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_byteenable;  // mm_interconnect_2:pll_stream_reconfig_mgmt_avalon_slave_byteenable -> pll_stream_reconfig:mgmt_byteenable
	wire          mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_write;       // mm_interconnect_2:pll_stream_reconfig_mgmt_avalon_slave_write -> pll_stream_reconfig:mgmt_write
	wire   [31:0] mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_writedata;   // mm_interconnect_2:pll_stream_reconfig_mgmt_avalon_slave_writedata -> pll_stream_reconfig:mgmt_writedata
	wire   [63:0] mm_interconnect_2_chip_id_read_mm_0_s0_readdata;                     // chip_id_read_mm_0:avs_s0_readdata -> mm_interconnect_2:chip_id_read_mm_0_s0_readdata
	wire          mm_interconnect_2_chip_id_read_mm_0_s0_read;                         // mm_interconnect_2:chip_id_read_mm_0_s0_read -> chip_id_read_mm_0:avs_s0_read
	wire   [31:0] mm_interconnect_2_hdmi_mm_bridge_s0_readdata;                        // hdmi_mm_bridge:s0_readdata -> mm_interconnect_2:hdmi_mm_bridge_s0_readdata
	wire          mm_interconnect_2_hdmi_mm_bridge_s0_waitrequest;                     // hdmi_mm_bridge:s0_waitrequest -> mm_interconnect_2:hdmi_mm_bridge_s0_waitrequest
	wire          mm_interconnect_2_hdmi_mm_bridge_s0_debugaccess;                     // mm_interconnect_2:hdmi_mm_bridge_s0_debugaccess -> hdmi_mm_bridge:s0_debugaccess
	wire   [12:0] mm_interconnect_2_hdmi_mm_bridge_s0_address;                         // mm_interconnect_2:hdmi_mm_bridge_s0_address -> hdmi_mm_bridge:s0_address
	wire          mm_interconnect_2_hdmi_mm_bridge_s0_read;                            // mm_interconnect_2:hdmi_mm_bridge_s0_read -> hdmi_mm_bridge:s0_read
	wire    [3:0] mm_interconnect_2_hdmi_mm_bridge_s0_byteenable;                      // mm_interconnect_2:hdmi_mm_bridge_s0_byteenable -> hdmi_mm_bridge:s0_byteenable
	wire          mm_interconnect_2_hdmi_mm_bridge_s0_readdatavalid;                   // hdmi_mm_bridge:s0_readdatavalid -> mm_interconnect_2:hdmi_mm_bridge_s0_readdatavalid
	wire          mm_interconnect_2_hdmi_mm_bridge_s0_write;                           // mm_interconnect_2:hdmi_mm_bridge_s0_write -> hdmi_mm_bridge:s0_write
	wire   [31:0] mm_interconnect_2_hdmi_mm_bridge_s0_writedata;                       // mm_interconnect_2:hdmi_mm_bridge_s0_writedata -> hdmi_mm_bridge:s0_writedata
	wire    [0:0] mm_interconnect_2_hdmi_mm_bridge_s0_burstcount;                      // mm_interconnect_2:hdmi_mm_bridge_s0_burstcount -> hdmi_mm_bridge:s0_burstcount
	wire          mm_interconnect_2_led_pio_s1_chipselect;                             // mm_interconnect_2:led_pio_s1_chipselect -> led_pio:chipselect
	wire   [31:0] mm_interconnect_2_led_pio_s1_readdata;                               // led_pio:readdata -> mm_interconnect_2:led_pio_s1_readdata
	wire    [1:0] mm_interconnect_2_led_pio_s1_address;                                // mm_interconnect_2:led_pio_s1_address -> led_pio:address
	wire          mm_interconnect_2_led_pio_s1_write;                                  // mm_interconnect_2:led_pio_s1_write -> led_pio:write_n
	wire   [31:0] mm_interconnect_2_led_pio_s1_writedata;                              // mm_interconnect_2:led_pio_s1_writedata -> led_pio:writedata
	wire          mm_interconnect_2_dipsw_pio_s1_chipselect;                           // mm_interconnect_2:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	wire   [31:0] mm_interconnect_2_dipsw_pio_s1_readdata;                             // dipsw_pio:readdata -> mm_interconnect_2:dipsw_pio_s1_readdata
	wire    [1:0] mm_interconnect_2_dipsw_pio_s1_address;                              // mm_interconnect_2:dipsw_pio_s1_address -> dipsw_pio:address
	wire          mm_interconnect_2_dipsw_pio_s1_write;                                // mm_interconnect_2:dipsw_pio_s1_write -> dipsw_pio:write_n
	wire   [31:0] mm_interconnect_2_dipsw_pio_s1_writedata;                            // mm_interconnect_2:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	wire          mm_interconnect_2_button_pio_s1_chipselect;                          // mm_interconnect_2:button_pio_s1_chipselect -> button_pio:chipselect
	wire   [31:0] mm_interconnect_2_button_pio_s1_readdata;                            // button_pio:readdata -> mm_interconnect_2:button_pio_s1_readdata
	wire    [1:0] mm_interconnect_2_button_pio_s1_address;                             // mm_interconnect_2:button_pio_s1_address -> button_pio:address
	wire          mm_interconnect_2_button_pio_s1_write;                               // mm_interconnect_2:button_pio_s1_write -> button_pio:write_n
	wire   [31:0] mm_interconnect_2_button_pio_s1_writedata;                           // mm_interconnect_2:button_pio_s1_writedata -> button_pio:writedata
	wire          mm_interconnect_2_pll_reset_pio_s1_chipselect;                       // mm_interconnect_2:pll_reset_pio_s1_chipselect -> pll_reset_pio:chipselect
	wire   [31:0] mm_interconnect_2_pll_reset_pio_s1_readdata;                         // pll_reset_pio:readdata -> mm_interconnect_2:pll_reset_pio_s1_readdata
	wire    [2:0] mm_interconnect_2_pll_reset_pio_s1_address;                          // mm_interconnect_2:pll_reset_pio_s1_address -> pll_reset_pio:address
	wire          mm_interconnect_2_pll_reset_pio_s1_write;                            // mm_interconnect_2:pll_reset_pio_s1_write -> pll_reset_pio:write_n
	wire   [31:0] mm_interconnect_2_pll_reset_pio_s1_writedata;                        // mm_interconnect_2:pll_reset_pio_s1_writedata -> pll_reset_pio:writedata
	wire          mm_interconnect_2_cvo_reset_pio_s1_chipselect;                       // mm_interconnect_2:cvo_reset_pio_s1_chipselect -> cvo_reset_pio:chipselect
	wire   [31:0] mm_interconnect_2_cvo_reset_pio_s1_readdata;                         // cvo_reset_pio:readdata -> mm_interconnect_2:cvo_reset_pio_s1_readdata
	wire    [2:0] mm_interconnect_2_cvo_reset_pio_s1_address;                          // mm_interconnect_2:cvo_reset_pio_s1_address -> cvo_reset_pio:address
	wire          mm_interconnect_2_cvo_reset_pio_s1_write;                            // mm_interconnect_2:cvo_reset_pio_s1_write -> cvo_reset_pio:write_n
	wire   [31:0] mm_interconnect_2_cvo_reset_pio_s1_writedata;                        // mm_interconnect_2:cvo_reset_pio_s1_writedata -> cvo_reset_pio:writedata
	wire   [31:0] mm_interconnect_2_locked_pio_s1_readdata;                            // locked_pio:readdata -> mm_interconnect_2:locked_pio_s1_readdata
	wire    [2:0] mm_interconnect_2_locked_pio_s1_address;                             // mm_interconnect_2:locked_pio_s1_address -> locked_pio:address
	wire          mm_interconnect_2_arduino_gpio_s1_chipselect;                        // mm_interconnect_2:arduino_gpio_s1_chipselect -> arduino_gpio:chipselect
	wire   [31:0] mm_interconnect_2_arduino_gpio_s1_readdata;                          // arduino_gpio:readdata -> mm_interconnect_2:arduino_gpio_s1_readdata
	wire    [2:0] mm_interconnect_2_arduino_gpio_s1_address;                           // mm_interconnect_2:arduino_gpio_s1_address -> arduino_gpio:address
	wire          mm_interconnect_2_arduino_gpio_s1_write;                             // mm_interconnect_2:arduino_gpio_s1_write -> arduino_gpio:write_n
	wire   [31:0] mm_interconnect_2_arduino_gpio_s1_writedata;                         // mm_interconnect_2:arduino_gpio_s1_writedata -> arduino_gpio:writedata
	wire          mm_interconnect_2_gpio_0_a_s1_chipselect;                            // mm_interconnect_2:gpio_0_a_s1_chipselect -> gpio_0_a:chipselect
	wire   [31:0] mm_interconnect_2_gpio_0_a_s1_readdata;                              // gpio_0_a:readdata -> mm_interconnect_2:gpio_0_a_s1_readdata
	wire    [2:0] mm_interconnect_2_gpio_0_a_s1_address;                               // mm_interconnect_2:gpio_0_a_s1_address -> gpio_0_a:address
	wire          mm_interconnect_2_gpio_0_a_s1_write;                                 // mm_interconnect_2:gpio_0_a_s1_write -> gpio_0_a:write_n
	wire   [31:0] mm_interconnect_2_gpio_0_a_s1_writedata;                             // mm_interconnect_2:gpio_0_a_s1_writedata -> gpio_0_a:writedata
	wire          mm_interconnect_2_gpio_0_b_s1_chipselect;                            // mm_interconnect_2:gpio_0_b_s1_chipselect -> gpio_0_b:chipselect
	wire   [31:0] mm_interconnect_2_gpio_0_b_s1_readdata;                              // gpio_0_b:readdata -> mm_interconnect_2:gpio_0_b_s1_readdata
	wire    [2:0] mm_interconnect_2_gpio_0_b_s1_address;                               // mm_interconnect_2:gpio_0_b_s1_address -> gpio_0_b:address
	wire          mm_interconnect_2_gpio_0_b_s1_write;                                 // mm_interconnect_2:gpio_0_b_s1_write -> gpio_0_b:write_n
	wire   [31:0] mm_interconnect_2_gpio_0_b_s1_writedata;                             // mm_interconnect_2:gpio_0_b_s1_writedata -> gpio_0_b:writedata
	wire          mm_interconnect_2_gpio_1_a_s1_chipselect;                            // mm_interconnect_2:gpio_1_a_s1_chipselect -> gpio_1_a:chipselect
	wire   [31:0] mm_interconnect_2_gpio_1_a_s1_readdata;                              // gpio_1_a:readdata -> mm_interconnect_2:gpio_1_a_s1_readdata
	wire    [2:0] mm_interconnect_2_gpio_1_a_s1_address;                               // mm_interconnect_2:gpio_1_a_s1_address -> gpio_1_a:address
	wire          mm_interconnect_2_gpio_1_a_s1_write;                                 // mm_interconnect_2:gpio_1_a_s1_write -> gpio_1_a:write_n
	wire   [31:0] mm_interconnect_2_gpio_1_a_s1_writedata;                             // mm_interconnect_2:gpio_1_a_s1_writedata -> gpio_1_a:writedata
	wire          mm_interconnect_2_gpio_1_b_s1_chipselect;                            // mm_interconnect_2:gpio_1_b_s1_chipselect -> gpio_1_b:chipselect
	wire   [31:0] mm_interconnect_2_gpio_1_b_s1_readdata;                              // gpio_1_b:readdata -> mm_interconnect_2:gpio_1_b_s1_readdata
	wire    [2:0] mm_interconnect_2_gpio_1_b_s1_address;                               // mm_interconnect_2:gpio_1_b_s1_address -> gpio_1_b:address
	wire          mm_interconnect_2_gpio_1_b_s1_write;                                 // mm_interconnect_2:gpio_1_b_s1_write -> gpio_1_b:write_n
	wire   [31:0] mm_interconnect_2_gpio_1_b_s1_writedata;                             // mm_interconnect_2:gpio_1_b_s1_writedata -> gpio_1_b:writedata
	wire          hdmi_mm_bridge_m0_waitrequest;                                       // mm_interconnect_3:hdmi_mm_bridge_m0_waitrequest -> hdmi_mm_bridge:m0_waitrequest
	wire   [31:0] hdmi_mm_bridge_m0_readdata;                                          // mm_interconnect_3:hdmi_mm_bridge_m0_readdata -> hdmi_mm_bridge:m0_readdata
	wire          hdmi_mm_bridge_m0_debugaccess;                                       // hdmi_mm_bridge:m0_debugaccess -> mm_interconnect_3:hdmi_mm_bridge_m0_debugaccess
	wire   [12:0] hdmi_mm_bridge_m0_address;                                           // hdmi_mm_bridge:m0_address -> mm_interconnect_3:hdmi_mm_bridge_m0_address
	wire          hdmi_mm_bridge_m0_read;                                              // hdmi_mm_bridge:m0_read -> mm_interconnect_3:hdmi_mm_bridge_m0_read
	wire    [3:0] hdmi_mm_bridge_m0_byteenable;                                        // hdmi_mm_bridge:m0_byteenable -> mm_interconnect_3:hdmi_mm_bridge_m0_byteenable
	wire          hdmi_mm_bridge_m0_readdatavalid;                                     // mm_interconnect_3:hdmi_mm_bridge_m0_readdatavalid -> hdmi_mm_bridge:m0_readdatavalid
	wire   [31:0] hdmi_mm_bridge_m0_writedata;                                         // hdmi_mm_bridge:m0_writedata -> mm_interconnect_3:hdmi_mm_bridge_m0_writedata
	wire          hdmi_mm_bridge_m0_write;                                             // hdmi_mm_bridge:m0_write -> mm_interconnect_3:hdmi_mm_bridge_m0_write
	wire    [0:0] hdmi_mm_bridge_m0_burstcount;                                        // hdmi_mm_bridge:m0_burstcount -> mm_interconnect_3:hdmi_mm_bridge_m0_burstcount
	wire   [31:0] mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_readdata;              // alt_vip_cl_vfb_hdmi:control_readdata -> mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_readdata
	wire          mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_waitrequest;           // alt_vip_cl_vfb_hdmi:control_waitrequest -> mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_waitrequest
	wire    [3:0] mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_address;               // mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_address -> alt_vip_cl_vfb_hdmi:control_address
	wire          mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_read;                  // mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_read -> alt_vip_cl_vfb_hdmi:control_read
	wire    [3:0] mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_byteenable;            // mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_byteenable -> alt_vip_cl_vfb_hdmi:control_byteenable
	wire          mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_readdatavalid;         // alt_vip_cl_vfb_hdmi:control_readdatavalid -> mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_readdatavalid
	wire          mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_write;                 // mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_write -> alt_vip_cl_vfb_hdmi:control_write
	wire   [31:0] mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_writedata;             // mm_interconnect_3:alt_vip_cl_vfb_hdmi_control_writedata -> alt_vip_cl_vfb_hdmi:control_writedata
	wire   [31:0] mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_readdata;              // alt_vip_cl_cvo_hdmi:control_readdata -> mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_readdata
	wire          mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_waitrequest;           // alt_vip_cl_cvo_hdmi:control_waitrequest -> mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_waitrequest
	wire    [7:0] mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_address;               // mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_address -> alt_vip_cl_cvo_hdmi:control_address
	wire          mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_read;                  // mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_read -> alt_vip_cl_cvo_hdmi:control_read
	wire    [3:0] mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_byteenable;            // mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_byteenable -> alt_vip_cl_cvo_hdmi:control_byteenable
	wire          mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_readdatavalid;         // alt_vip_cl_cvo_hdmi:control_readdatavalid -> mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_readdatavalid
	wire          mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_write;                 // mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_write -> alt_vip_cl_cvo_hdmi:control_write
	wire   [31:0] mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_writedata;             // mm_interconnect_3:alt_vip_cl_cvo_hdmi_control_writedata -> alt_vip_cl_cvo_hdmi:control_writedata
	wire          custom_ip_bridge_m0_waitrequest;                                     // mm_interconnect_4:custom_ip_bridge_m0_waitrequest -> custom_ip_bridge:m0_waitrequest
	wire   [31:0] custom_ip_bridge_m0_readdata;                                        // mm_interconnect_4:custom_ip_bridge_m0_readdata -> custom_ip_bridge:m0_readdata
	wire          custom_ip_bridge_m0_debugaccess;                                     // custom_ip_bridge:m0_debugaccess -> mm_interconnect_4:custom_ip_bridge_m0_debugaccess
	wire    [5:0] custom_ip_bridge_m0_address;                                         // custom_ip_bridge:m0_address -> mm_interconnect_4:custom_ip_bridge_m0_address
	wire          custom_ip_bridge_m0_read;                                            // custom_ip_bridge:m0_read -> mm_interconnect_4:custom_ip_bridge_m0_read
	wire    [3:0] custom_ip_bridge_m0_byteenable;                                      // custom_ip_bridge:m0_byteenable -> mm_interconnect_4:custom_ip_bridge_m0_byteenable
	wire          custom_ip_bridge_m0_readdatavalid;                                   // mm_interconnect_4:custom_ip_bridge_m0_readdatavalid -> custom_ip_bridge:m0_readdatavalid
	wire   [31:0] custom_ip_bridge_m0_writedata;                                       // custom_ip_bridge:m0_writedata -> mm_interconnect_4:custom_ip_bridge_m0_writedata
	wire          custom_ip_bridge_m0_write;                                           // custom_ip_bridge:m0_write -> mm_interconnect_4:custom_ip_bridge_m0_write
	wire    [0:0] custom_ip_bridge_m0_burstcount;                                      // custom_ip_bridge:m0_burstcount -> mm_interconnect_4:custom_ip_bridge_m0_burstcount
	wire   [31:0] mm_interconnect_4_random_s1_readdata;                                // random:readdata -> mm_interconnect_4:random_s1_readdata
	wire    [1:0] mm_interconnect_4_random_s1_address;                                 // mm_interconnect_4:random_s1_address -> random:address
	wire          mm_interconnect_4_ctrl_register_s1_chipselect;                       // mm_interconnect_4:ctrl_register_s1_chipselect -> ctrl_register:chipselect
	wire   [31:0] mm_interconnect_4_ctrl_register_s1_readdata;                         // ctrl_register:readdata -> mm_interconnect_4:ctrl_register_s1_readdata
	wire    [1:0] mm_interconnect_4_ctrl_register_s1_address;                          // mm_interconnect_4:ctrl_register_s1_address -> ctrl_register:address
	wire          mm_interconnect_4_ctrl_register_s1_write;                            // mm_interconnect_4:ctrl_register_s1_write -> ctrl_register:write_n
	wire   [31:0] mm_interconnect_4_ctrl_register_s1_writedata;                        // mm_interconnect_4:ctrl_register_s1_writedata -> ctrl_register:writedata
	wire          mm_interconnect_4_lfsr_reset_value_reg_s1_chipselect;                // mm_interconnect_4:lfsr_reset_value_reg_s1_chipselect -> lfsr_reset_value_reg:chipselect
	wire   [31:0] mm_interconnect_4_lfsr_reset_value_reg_s1_readdata;                  // lfsr_reset_value_reg:readdata -> mm_interconnect_4:lfsr_reset_value_reg_s1_readdata
	wire    [1:0] mm_interconnect_4_lfsr_reset_value_reg_s1_address;                   // mm_interconnect_4:lfsr_reset_value_reg_s1_address -> lfsr_reset_value_reg:address
	wire          mm_interconnect_4_lfsr_reset_value_reg_s1_write;                     // mm_interconnect_4:lfsr_reset_value_reg_s1_write -> lfsr_reset_value_reg:write_n
	wire   [31:0] mm_interconnect_4_lfsr_reset_value_reg_s1_writedata;                 // mm_interconnect_4:lfsr_reset_value_reg_s1_writedata -> lfsr_reset_value_reg:writedata
	wire          alt_vip_cl_vfb_hdmi_mem_master_rd_waitrequest;                       // mm_interconnect_5:alt_vip_cl_vfb_hdmi_mem_master_rd_waitrequest -> alt_vip_cl_vfb_hdmi:mem_master_rd_waitrequest
	wire  [255:0] alt_vip_cl_vfb_hdmi_mem_master_rd_readdata;                          // mm_interconnect_5:alt_vip_cl_vfb_hdmi_mem_master_rd_readdata -> alt_vip_cl_vfb_hdmi:mem_master_rd_readdata
	wire   [31:0] alt_vip_cl_vfb_hdmi_mem_master_rd_address;                           // alt_vip_cl_vfb_hdmi:mem_master_rd_address -> mm_interconnect_5:alt_vip_cl_vfb_hdmi_mem_master_rd_address
	wire          alt_vip_cl_vfb_hdmi_mem_master_rd_read;                              // alt_vip_cl_vfb_hdmi:mem_master_rd_read -> mm_interconnect_5:alt_vip_cl_vfb_hdmi_mem_master_rd_read
	wire          alt_vip_cl_vfb_hdmi_mem_master_rd_readdatavalid;                     // mm_interconnect_5:alt_vip_cl_vfb_hdmi_mem_master_rd_readdatavalid -> alt_vip_cl_vfb_hdmi:mem_master_rd_readdatavalid
	wire    [5:0] alt_vip_cl_vfb_hdmi_mem_master_rd_burstcount;                        // alt_vip_cl_vfb_hdmi:mem_master_rd_burstcount -> mm_interconnect_5:alt_vip_cl_vfb_hdmi_mem_master_rd_burstcount
	wire  [255:0] mm_interconnect_5_hps_0_f2h_sdram0_data_readdata;                    // hps_0:f2h_sdram0_READDATA -> mm_interconnect_5:hps_0_f2h_sdram0_data_readdata
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_waitrequest;                 // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_5:hps_0_f2h_sdram0_data_waitrequest
	wire   [26:0] mm_interconnect_5_hps_0_f2h_sdram0_data_address;                     // mm_interconnect_5:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_read;                        // mm_interconnect_5:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	wire   [31:0] mm_interconnect_5_hps_0_f2h_sdram0_data_byteenable;                  // mm_interconnect_5:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_readdatavalid;               // hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_5:hps_0_f2h_sdram0_data_readdatavalid
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_write;                       // mm_interconnect_5:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire  [255:0] mm_interconnect_5_hps_0_f2h_sdram0_data_writedata;                   // mm_interconnect_5:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_burstcount;                  // mm_interconnect_5:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire          irq_mapper_receiver0_irq;                                            // alt_vip_cl_vfb_hdmi:control_interrupt_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                            // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                            // dipsw_pio:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                            // button_pio:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                            // arduino_gpio:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                            // alt_vip_cl_cvo_hdmi:status_update_irq_irq -> irq_mapper:receiver5_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                                  // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                  // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          altchip_id_0_output_valid;                                           // altchip_id_0:data_valid -> avalon_st_adapter:in_0_valid
	wire   [63:0] altchip_id_0_output_data;                                            // altchip_id_0:chip_id -> avalon_st_adapter:in_0_data
	wire   [63:0] avalon_st_adapter_out_0_data;                                        // avalon_st_adapter:out_0_data -> chip_id_read_mm_0:asi_in0_data
	wire          avalon_st_adapter_out_0_ready;                                       // chip_id_read_mm_0:asi_in0_ready -> avalon_st_adapter:out_0_ready
	wire          rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [alt_vip_cl_vfb_hdmi:mem_reset, mm_interconnect_5:alt_vip_cl_vfb_hdmi_mem_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [altchip_id_0:reset, arduino_gpio:reset_n, avalon_st_adapter:in_rst_0_reset, button_pio:reset_n, chip_id_read_mm_0:reset, ctrl_register:reset_n, custom_ip_bridge:reset, cvo_reset_pio:reset_n, dipsw_pio:reset_n, gpio_0_a:reset_n, gpio_0_b:reset_n, gpio_1_a:reset_n, gpio_1_b:reset_n, jtag_uart:rst_n, led_pio:reset_n, lfsr_reset_value_reg:reset_n, locked_pio:reset_n, lw_mm_bridge:reset, mm_interconnect_0:custom_ip_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:lw_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_2:lw_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_4:custom_ip_bridge_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, pll_reset_pio:reset_n, pll_stream_reconfig:mgmt_reset, random:reset_n, rst_translator:in_reset, sysid_qsys:reset_n]
	wire          rst_controller_001_reset_out_reset_req;                              // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_002_reset_out_reset;                                  // rst_controller_002:reset_out -> [rst_controller_001:reset_in0, rst_controller_003:reset_in0]
	wire          hps_0_h2f_reset_reset;                                               // hps_0:h2f_rst_n -> [rst_controller_002:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0]
	wire          por_reset_reset;                                                     // por:reset -> rst_controller_002:reset_in1
	wire          rst_controller_003_reset_out_reset;                                  // rst_controller_003:reset_out -> custom_reset_synchronizer:reset_in
	wire          rst_controller_004_reset_out_reset;                                  // rst_controller_004:reset_out -> rst_controller_004_reset_out_reset:in
	wire          rst_controller_005_reset_out_reset;                                  // rst_controller_005:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_006_reset_out_reset;                                  // rst_controller_006:reset_out -> mm_interconnect_5:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset

	soc_system_alt_vip_cl_cvo_hdmi #(
		.BPS                           (8),
		.NUMBER_OF_COLOUR_PLANES       (4),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1920),
		.V_ACTIVE_LINES                (1080),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (1920),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (1),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (1919),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.ACCEPT_SYNC                   (0),
		.COUNT_STEP_IS_PIP_VALUE       (0),
		.LOW_LATENCY                   (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (32),
		.H_FRONT_PORCH                 (32),
		.H_BACK_PORCH                  (64),
		.V_SYNC_LENGTH                 (3),
		.V_FRONT_PORCH                 (1),
		.V_BACK_PORCH                  (27),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0),
		.PIXELS_IN_PARALLEL            (1),
		.SRC_WIDTH                     (8),
		.DST_WIDTH                     (8),
		.CONTEXT_WIDTH                 (8),
		.TASK_WIDTH                    (8)
	) alt_vip_cl_cvo_hdmi (
		.clocked_video_vid_clk         (alt_vip_cl_cvo_hdmi_clocked_video_vid_clk),                   //     clocked_video.vid_clk
		.clocked_video_vid_data        (alt_vip_cl_cvo_hdmi_clocked_video_vid_data),                  //                  .vid_data
		.clocked_video_underflow       (alt_vip_cl_cvo_hdmi_clocked_video_underflow),                 //                  .underflow
		.clocked_video_vid_mode_change (alt_vip_cl_cvo_hdmi_clocked_video_vid_mode_change),           //                  .vid_mode_change
		.clocked_video_vid_std         (alt_vip_cl_cvo_hdmi_clocked_video_vid_std),                   //                  .vid_std
		.clocked_video_vid_datavalid   (alt_vip_cl_cvo_hdmi_clocked_video_vid_datavalid),             //                  .vid_datavalid
		.clocked_video_vid_v_sync      (alt_vip_cl_cvo_hdmi_clocked_video_vid_v_sync),                //                  .vid_v_sync
		.clocked_video_vid_h_sync      (alt_vip_cl_cvo_hdmi_clocked_video_vid_h_sync),                //                  .vid_h_sync
		.clocked_video_vid_f           (alt_vip_cl_cvo_hdmi_clocked_video_vid_f),                     //                  .vid_f
		.clocked_video_vid_h           (alt_vip_cl_cvo_hdmi_clocked_video_vid_h),                     //                  .vid_h
		.clocked_video_vid_v           (alt_vip_cl_cvo_hdmi_clocked_video_vid_v),                     //                  .vid_v
		.main_clock_clk                (clk_hdmi_clk),                                                //        main_clock.clk
		.main_reset_reset              (custom_reset_synchronizer_reset_out_reset),                   //        main_reset.reset
		.din_data                      (alt_vip_cl_vfb_hdmi_dout_data),                               //               din.data
		.din_valid                     (alt_vip_cl_vfb_hdmi_dout_valid),                              //                  .valid
		.din_startofpacket             (alt_vip_cl_vfb_hdmi_dout_startofpacket),                      //                  .startofpacket
		.din_endofpacket               (alt_vip_cl_vfb_hdmi_dout_endofpacket),                        //                  .endofpacket
		.din_ready                     (alt_vip_cl_vfb_hdmi_dout_ready),                              //                  .ready
		.control_address               (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_address),       //           control.address
		.control_byteenable            (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_byteenable),    //                  .byteenable
		.control_write                 (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_write),         //                  .write
		.control_writedata             (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_writedata),     //                  .writedata
		.control_read                  (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_read),          //                  .read
		.control_readdata              (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_readdata),      //                  .readdata
		.control_readdatavalid         (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_readdatavalid), //                  .readdatavalid
		.control_waitrequest           (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_waitrequest),   //                  .waitrequest
		.status_update_irq_irq         (irq_mapper_receiver5_irq)                                     // status_update_irq.irq
	);

	soc_system_alt_vip_cl_vfb_hdmi #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (4),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.READY_LATENCY                (1),
		.MAX_WIDTH                    (1920),
		.MAX_HEIGHT                   (1080),
		.CLOCKS_ARE_SEPARATE          (1),
		.MEM_PORT_WIDTH               (256),
		.MEM_BASE_ADDR                (0),
		.BURST_ALIGNMENT              (1),
		.WRITE_FIFO_DEPTH             (8),
		.WRITE_BURST_TARGET           (2),
		.READ_FIFO_DEPTH              (256),
		.READ_BURST_TARGET            (32),
		.WRITER_RUNTIME_CONTROL       (0),
		.READER_RUNTIME_CONTROL       (1),
		.IS_FRAME_WRITER              (0),
		.IS_FRAME_READER              (1),
		.DROP_FRAMES                  (0),
		.REPEAT_FRAMES                (1),
		.DROP_REPEAT_USER             (0),
		.INTERLACED_SUPPORT           (0),
		.CONTROLLED_DROP_REPEAT       (0),
		.DROP_INVALID_FIELDS          (0),
		.MULTI_FRAME_DELAY            (1),
		.IS_SYNC_MASTER               (0),
		.IS_SYNC_SLAVE                (0),
		.LINE_BASED_BUFFERING         (0),
		.PRIORITIZE_FMAX              (0),
		.USER_PACKETS_MAX_STORAGE     (0),
		.MAX_SYMBOLS_PER_PACKET       (10),
		.NUM_BUFFERS                  (3)
	) alt_vip_cl_vfb_hdmi (
		.main_clock                  (clk_hdmi_clk),                                                //        main_clock.clk
		.main_reset                  (custom_reset_synchronizer_reset_out_reset),                   //        main_reset.reset
		.mem_clock                   (hps_0_h2f_user0_clock_clk),                                   //         mem_clock.clk
		.mem_reset                   (rst_controller_reset_out_reset),                              //         mem_reset.reset
		.dout_data                   (alt_vip_cl_vfb_hdmi_dout_data),                               //              dout.data
		.dout_valid                  (alt_vip_cl_vfb_hdmi_dout_valid),                              //                  .valid
		.dout_startofpacket          (alt_vip_cl_vfb_hdmi_dout_startofpacket),                      //                  .startofpacket
		.dout_endofpacket            (alt_vip_cl_vfb_hdmi_dout_endofpacket),                        //                  .endofpacket
		.dout_ready                  (alt_vip_cl_vfb_hdmi_dout_ready),                              //                  .ready
		.mem_master_rd_address       (alt_vip_cl_vfb_hdmi_mem_master_rd_address),                   //     mem_master_rd.address
		.mem_master_rd_burstcount    (alt_vip_cl_vfb_hdmi_mem_master_rd_burstcount),                //                  .burstcount
		.mem_master_rd_waitrequest   (alt_vip_cl_vfb_hdmi_mem_master_rd_waitrequest),               //                  .waitrequest
		.mem_master_rd_read          (alt_vip_cl_vfb_hdmi_mem_master_rd_read),                      //                  .read
		.mem_master_rd_readdata      (alt_vip_cl_vfb_hdmi_mem_master_rd_readdata),                  //                  .readdata
		.mem_master_rd_readdatavalid (alt_vip_cl_vfb_hdmi_mem_master_rd_readdatavalid),             //                  .readdatavalid
		.control_interrupt_irq       (irq_mapper_receiver0_irq),                                    // control_interrupt.irq
		.control_address             (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_address),       //           control.address
		.control_byteenable          (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_byteenable),    //                  .byteenable
		.control_write               (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_write),         //                  .write
		.control_writedata           (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_writedata),     //                  .writedata
		.control_read                (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_read),          //                  .read
		.control_readdata            (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_readdata),      //                  .readdata
		.control_readdatavalid       (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_readdatavalid), //                  .readdatavalid
		.control_waitrequest         (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_waitrequest)    //                  .waitrequest
	);

	altchip_id #(
		.DEVICE_FAMILY ("Cyclone V"),
		.ID_VALUE      (64'b1111111111111111111111111111111111111111111111111111111111111111)
	) altchip_id_0 (
		.clkin      (clk_clk),                            //  clkin.clk
		.reset      (rst_controller_001_reset_out_reset), //  reset.reset
		.data_valid (altchip_id_0_output_valid),          // output.valid
		.chip_id    (altchip_id_0_output_data)            //       .data
	);

	soc_system_arduino_gpio arduino_gpio (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_2_arduino_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_arduino_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_arduino_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_arduino_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_arduino_gpio_s1_readdata),   //                    .readdata
		.bidir_port (arduino_gpio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                      //                 irq.irq
	);

	soc_system_button_pio button_pio (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_2_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                    //                 irq.irq
	);

	chip_id_read_mm chip_id_read_mm_0 (
		.clk             (clk_clk),                                         // clock.clk
		.reset           (rst_controller_001_reset_out_reset),              // reset.reset
		.avs_s0_read     (mm_interconnect_2_chip_id_read_mm_0_s0_read),     //    s0.read
		.avs_s0_readdata (mm_interconnect_2_chip_id_read_mm_0_s0_readdata), //      .readdata
		.asi_in0_data    (avalon_st_adapter_out_0_data),                    //   in0.data
		.asi_in0_ready   (avalon_st_adapter_out_0_ready)                    //      .ready
	);

	soc_system_ctrl_register ctrl_register (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_4_ctrl_register_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_4_ctrl_register_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_4_ctrl_register_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_4_ctrl_register_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_4_ctrl_register_s1_readdata),   //                    .readdata
		.out_port   (ctrl_reg_export)                                // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (6),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) custom_ip_bridge (
		.clk              (clk_clk),                                             //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_0_custom_ip_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_custom_ip_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_custom_ip_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_custom_ip_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_custom_ip_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_custom_ip_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_custom_ip_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_custom_ip_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_custom_ip_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_custom_ip_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (custom_ip_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (custom_ip_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (custom_ip_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (custom_ip_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (custom_ip_bridge_m0_writedata),                       //      .writedata
		.m0_address       (custom_ip_bridge_m0_address),                         //      .address
		.m0_write         (custom_ip_bridge_m0_write),                           //      .write
		.m0_read          (custom_ip_bridge_m0_read),                            //      .read
		.m0_byteenable    (custom_ip_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (custom_ip_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                    // (terminated)
		.m0_response      (2'b00)                                                // (terminated)
	);

	reset_sync_block #(
		.SYNC_DEPTH             (3),
		.ADDITIONAL_DEPTH       (2),
		.DISABLE_GLOBAL_NETWORK (1),
		.SYNC_BOTH_EDGES        (0)
	) custom_reset_synchronizer (
		.clk_in    (pll_stream_outclk0_clk),                    //  clock_in.clk
		.reset_in  (rst_controller_003_reset_out_reset),        //  reset_in.reset
		.clk_out   (clk_hdmi_clk),                              // clock_out.clk
		.reset_out (custom_reset_synchronizer_reset_out_reset)  // reset_out.reset
	);

	soc_system_cvo_reset_pio cvo_reset_pio (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_2_cvo_reset_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_cvo_reset_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_cvo_reset_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_cvo_reset_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_cvo_reset_pio_s1_readdata),   //                    .readdata
		.out_port   (cvo_reset_pio_external_connection_export)       // external_connection.export
	);

	soc_system_dipsw_pio dipsw_pio (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_2_dipsw_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_dipsw_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_dipsw_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_dipsw_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_dipsw_pio_s1_readdata),   //                    .readdata
		.in_port    (dipsw_pio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	soc_system_gpio_0_a gpio_0_a (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_gpio_0_a_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_gpio_0_a_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_gpio_0_a_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_gpio_0_a_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_gpio_0_a_s1_readdata),   //                    .readdata
		.bidir_port (gpio_0_a_export)                           // external_connection.export
	);

	soc_system_gpio_0_a gpio_0_b (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_gpio_0_b_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_gpio_0_b_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_gpio_0_b_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_gpio_0_b_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_gpio_0_b_s1_readdata),   //                    .readdata
		.bidir_port (gpio_0_b_export)                           // external_connection.export
	);

	soc_system_gpio_0_a gpio_1_a (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_gpio_1_a_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_gpio_1_a_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_gpio_1_a_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_gpio_1_a_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_gpio_1_a_s1_readdata),   //                    .readdata
		.bidir_port (gpio_1_a_export)                           // external_connection.export
	);

	soc_system_gpio_0_a gpio_1_b (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_gpio_1_b_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_gpio_1_b_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_gpio_1_b_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_gpio_1_b_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_gpio_1_b_s1_readdata),   //                    .readdata
		.bidir_port (gpio_1_b_export)                           // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (13),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) hdmi_mm_bridge (
		.clk              (clk_hdmi_clk),                                      //   clk.clk
		.reset            (custom_reset_synchronizer_reset_out_reset),         // reset.reset
		.s0_waitrequest   (mm_interconnect_2_hdmi_mm_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_2_hdmi_mm_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_2_hdmi_mm_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_2_hdmi_mm_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_2_hdmi_mm_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_2_hdmi_mm_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_2_hdmi_mm_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_2_hdmi_mm_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_2_hdmi_mm_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_2_hdmi_mm_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (hdmi_mm_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (hdmi_mm_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (hdmi_mm_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (hdmi_mm_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (hdmi_mm_bridge_m0_writedata),                       //      .writedata
		.m0_address       (hdmi_mm_bridge_m0_address),                         //      .address
		.m0_write         (hdmi_mm_bridge_m0_write),                           //      .write
		.m0_read          (hdmi_mm_bridge_m0_read),                            //      .read
		.m0_byteenable    (hdmi_mm_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (hdmi_mm_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                  // (terminated)
		.m0_response      (2'b00)                                              // (terminated)
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),                      //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),                     // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),                      //  f2h_warm_reset_req.reset_n
		.h2f_user0_clk            (hps_0_h2f_user0_clock_clk),                             //     h2f_user0_clock.clk
		.h2f_user1_clk            (hps_0_h2f_user1_clock_clk),                             //     h2f_user1_clock.clk
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),                  //   f2h_stm_hw_events.stm_hwevents
		.spim0_txd                (hps_0_spim0_txd),                                       //               spim0.txd
		.spim0_rxd                (hps_0_spim0_rxd),                                       //                    .rxd
		.spim0_ss_in_n            (hps_0_spim0_ss_in_n),                                   //                    .ss_in_n
		.spim0_ssi_oe_n           (hps_0_spim0_ssi_oe_n),                                  //                    .ssi_oe_n
		.spim0_ss_0_n             (hps_0_spim0_ss_0_n),                                    //                    .ss_0_n
		.spim0_ss_1_n             (hps_0_spim0_ss_1_n),                                    //                    .ss_1_n
		.spim0_ss_2_n             (hps_0_spim0_ss_2_n),                                    //                    .ss_2_n
		.spim0_ss_3_n             (hps_0_spim0_ss_3_n),                                    //                    .ss_3_n
		.spim0_sclk_out           (hps_0_spim0_sclk_out_clk),                              //      spim0_sclk_out.clk
		.uart1_cts                (hps_0_uart1_cts),                                       //               uart1.cts
		.uart1_dsr                (hps_0_uart1_dsr),                                       //                    .dsr
		.uart1_dcd                (hps_0_uart1_dcd),                                       //                    .dcd
		.uart1_ri                 (hps_0_uart1_ri),                                        //                    .ri
		.uart1_dtr                (hps_0_uart1_dtr),                                       //                    .dtr
		.uart1_rts                (hps_0_uart1_rts),                                       //                    .rts
		.uart1_out1_n             (hps_0_uart1_out1_n),                                    //                    .out1_n
		.uart1_out2_n             (hps_0_uart1_out2_n),                                    //                    .out2_n
		.uart1_rxd                (hps_0_uart1_rxd),                                       //                    .rxd
		.uart1_txd                (hps_0_uart1_txd),                                       //                    .txd
		.i2c_emac0_scl            (hps_0_i2c2_scl_in_clk),                                 //         i2c2_scl_in.clk
		.i2c_emac0_out_clk        (hps_0_i2c2_clk_clk),                                    //            i2c2_clk.clk
		.i2c_emac0_out_data       (hps_0_i2c2_out_data),                                   //                i2c2.out_data
		.i2c_emac0_sda            (hps_0_i2c2_sda),                                        //                    .sda
		.i2c_emac1_scl            (hps_0_i2c3_scl_in_clk),                                 //         i2c3_scl_in.clk
		.i2c_emac1_out_clk        (hps_0_i2c3_clk_clk),                                    //            i2c3_clk.clk
		.i2c_emac1_out_data       (hps_0_i2c3_out_data),                                   //                i2c3.out_data
		.i2c_emac1_sda            (hps_0_i2c3_sda),                                        //                    .sda
		.mem_a                    (memory_mem_a),                                          //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                         //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                         //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                       //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                        //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                       //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                      //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                      //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                       //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                    //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                         //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                        //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                      //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                        //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                         //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                      //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),                 //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),                   //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),                   //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),                   //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),                   //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),                   //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),                   //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),                    //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),                 //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),                 //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),                 //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),                   //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),                   //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),                   //                    .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),                     //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),                      //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),                      //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),                     //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),                      //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),                      //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),                      //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),                      //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),                      //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),                      //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),                      //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),                      //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),                      //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),                      //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),                     //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),                     //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),                     //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),                     //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),                    //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),                   //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),                   //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),                    //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),                     //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),                     //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),                     //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),                     //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),                     //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),                     //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),                  //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                  //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),                  //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                  //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                  //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),                  //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),                                 //           h2f_reset.reset_n
		.f2h_sdram0_clk           (hps_0_h2f_user0_clock_clk),                             //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_5_hps_0_f2h_sdram0_data_address),       //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_5_hps_0_f2h_sdram0_data_burstcount),    //                    .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_5_hps_0_f2h_sdram0_data_waitrequest),   //                    .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_5_hps_0_f2h_sdram0_data_readdata),      //                    .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_5_hps_0_f2h_sdram0_data_readdatavalid), //                    .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_5_hps_0_f2h_sdram0_data_read),          //                    .read
		.f2h_sdram0_WRITEDATA     (mm_interconnect_5_hps_0_f2h_sdram0_data_writedata),     //                    .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_5_hps_0_f2h_sdram0_data_byteenable),    //                    .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_5_hps_0_f2h_sdram0_data_write),         //                    .write
		.h2f_axi_clk              (clk_clk),                                               //       h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                             //      h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                           //                    .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                            //                    .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                           //                    .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                          //                    .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                           //                    .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                          //                    .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                           //                    .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                          //                    .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                          //                    .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                              //                    .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                            //                    .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                            //                    .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                            //                    .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                           //                    .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                           //                    .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                              //                    .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                            //                    .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                           //                    .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                           //                    .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                             //                    .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                           //                    .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                            //                    .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                           //                    .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                          //                    .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                           //                    .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                          //                    .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                           //                    .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                          //                    .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                          //                    .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                              //                    .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                            //                    .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                            //                    .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                            //                    .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                           //                    .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                           //                    .rready
		.f2h_axi_clk              (hps_0_h2f_user0_clock_clk),                             //       f2h_axi_clock.clk
		.f2h_AWID                 (),                                                      //       f2h_axi_slave.awid
		.f2h_AWADDR               (),                                                      //                    .awaddr
		.f2h_AWLEN                (),                                                      //                    .awlen
		.f2h_AWSIZE               (),                                                      //                    .awsize
		.f2h_AWBURST              (),                                                      //                    .awburst
		.f2h_AWLOCK               (),                                                      //                    .awlock
		.f2h_AWCACHE              (),                                                      //                    .awcache
		.f2h_AWPROT               (),                                                      //                    .awprot
		.f2h_AWVALID              (),                                                      //                    .awvalid
		.f2h_AWREADY              (),                                                      //                    .awready
		.f2h_AWUSER               (),                                                      //                    .awuser
		.f2h_WID                  (),                                                      //                    .wid
		.f2h_WDATA                (),                                                      //                    .wdata
		.f2h_WSTRB                (),                                                      //                    .wstrb
		.f2h_WLAST                (),                                                      //                    .wlast
		.f2h_WVALID               (),                                                      //                    .wvalid
		.f2h_WREADY               (),                                                      //                    .wready
		.f2h_BID                  (),                                                      //                    .bid
		.f2h_BRESP                (),                                                      //                    .bresp
		.f2h_BVALID               (),                                                      //                    .bvalid
		.f2h_BREADY               (),                                                      //                    .bready
		.f2h_ARID                 (),                                                      //                    .arid
		.f2h_ARADDR               (),                                                      //                    .araddr
		.f2h_ARLEN                (),                                                      //                    .arlen
		.f2h_ARSIZE               (),                                                      //                    .arsize
		.f2h_ARBURST              (),                                                      //                    .arburst
		.f2h_ARLOCK               (),                                                      //                    .arlock
		.f2h_ARCACHE              (),                                                      //                    .arcache
		.f2h_ARPROT               (),                                                      //                    .arprot
		.f2h_ARVALID              (),                                                      //                    .arvalid
		.f2h_ARREADY              (),                                                      //                    .arready
		.f2h_ARUSER               (),                                                      //                    .aruser
		.f2h_RID                  (),                                                      //                    .rid
		.f2h_RDATA                (),                                                      //                    .rdata
		.f2h_RRESP                (),                                                      //                    .rresp
		.f2h_RLAST                (),                                                      //                    .rlast
		.f2h_RVALID               (),                                                      //                    .rvalid
		.f2h_RREADY               (),                                                      //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                                               //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                          //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                        //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                         //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                        //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                       //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                        //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                       //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                        //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                       //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                       //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                           //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                         //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                         //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                         //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                        //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                        //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                           //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                         //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                        //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                        //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                          //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                        //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                         //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                        //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                       //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                        //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                       //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                        //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                       //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                       //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                           //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                         //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                         //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                         //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                        //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                        //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                                    //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                                     //            f2h_irq1.irq
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_2_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_2_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_2_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_2_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_2_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_2_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_2_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	soc_system_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_2_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	soc_system_lfsr_reset_value_reg lfsr_reset_value_reg (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_4_lfsr_reset_value_reg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_4_lfsr_reset_value_reg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_4_lfsr_reset_value_reg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_4_lfsr_reset_value_reg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_4_lfsr_reset_value_reg_s1_readdata),   //                    .readdata
		.out_port   (reset_val_export)                                      // external_connection.export
	);

	soc_system_locked_pio locked_pio (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_2_locked_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_locked_pio_s1_readdata), //                    .readdata
		.in_port  (pll_stream_locked_export)                  // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (17),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) lw_mm_bridge (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),              // reset.reset
		.s0_waitrequest   (mm_interconnect_1_lw_mm_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_lw_mm_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_lw_mm_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_lw_mm_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_lw_mm_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_lw_mm_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_lw_mm_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_lw_mm_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_lw_mm_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_lw_mm_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (lw_mm_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (lw_mm_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (lw_mm_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (lw_mm_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (lw_mm_bridge_m0_writedata),                       //      .writedata
		.m0_address       (lw_mm_bridge_m0_address),                         //      .address
		.m0_write         (lw_mm_bridge_m0_write),                           //      .write
		.m0_read          (lw_mm_bridge_m0_read),                            //      .read
		.m0_byteenable    (lw_mm_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (lw_mm_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                // (terminated)
		.m0_response      (2'b00)                                            // (terminated)
	);

	soc_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	soc_system_cvo_reset_pio pll_reset_pio (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_2_pll_reset_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_pll_reset_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_pll_reset_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_pll_reset_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_pll_reset_pio_s1_readdata),   //                    .readdata
		.out_port   (pll_reset_pio_external_connection_export)       // external_connection.export
	);

	soc_system_pll_stream pll_stream (
		.refclk            (clk_clk),                                             //            refclk.clk
		.rst               (pll_reset_pio_external_connection_export),            //             reset.reset
		.outclk_0          (pll_stream_outclk0_clk),                              //           outclk0.clk
		.locked            (pll_stream_locked_export),                            //            locked.export
		.reconfig_to_pll   (pll_stream_reconfig_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_stream_reconfig_from_pll_reconfig_from_pll)       // reconfig_from_pll.reconfig_from_pll
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (1),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_stream_reconfig (
		.mgmt_clk          (clk_clk),                                                             //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_001_reset_out_reset),                                  //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_writedata),   //                  .writedata
		.mgmt_byteenable   (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_byteenable),  //                  .byteenable
		.reconfig_to_pll   (pll_stream_reconfig_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_stream_reconfig_from_pll_reconfig_from_pll)                       // reconfig_from_pll.reconfig_from_pll
	);

	power_on_reset #(
		.POR_COUNT (20)
	) por (
		.clk   (clk_clk),         // clock.clk
		.reset (por_reset_reset)  // reset.reset
	);

	soc_system_random random (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_4_random_s1_address),  //                  s1.address
		.readdata (mm_interconnect_4_random_s1_readdata), //                    .readdata
		.in_port  (random_reg_export)                     // external_connection.export
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                           //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                         //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                          //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                         //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                        //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                         //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                        //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                         //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                        //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                        //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                            //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                          //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                          //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                          //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                         //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                         //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                            //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                          //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                         //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                         //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                           //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                         //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                          //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                         //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                        //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                         //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                        //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                         //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                        //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                        //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                            //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                          //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                          //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                          //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                         //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                         //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                             //                                                  clk_0_clk.clk
		.custom_ip_bridge_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                  //               custom_ip_bridge_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                  // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.custom_ip_bridge_s0_address                                      (mm_interconnect_0_custom_ip_bridge_s0_address),       //                                        custom_ip_bridge_s0.address
		.custom_ip_bridge_s0_write                                        (mm_interconnect_0_custom_ip_bridge_s0_write),         //                                                           .write
		.custom_ip_bridge_s0_read                                         (mm_interconnect_0_custom_ip_bridge_s0_read),          //                                                           .read
		.custom_ip_bridge_s0_readdata                                     (mm_interconnect_0_custom_ip_bridge_s0_readdata),      //                                                           .readdata
		.custom_ip_bridge_s0_writedata                                    (mm_interconnect_0_custom_ip_bridge_s0_writedata),     //                                                           .writedata
		.custom_ip_bridge_s0_burstcount                                   (mm_interconnect_0_custom_ip_bridge_s0_burstcount),    //                                                           .burstcount
		.custom_ip_bridge_s0_byteenable                                   (mm_interconnect_0_custom_ip_bridge_s0_byteenable),    //                                                           .byteenable
		.custom_ip_bridge_s0_readdatavalid                                (mm_interconnect_0_custom_ip_bridge_s0_readdatavalid), //                                                           .readdatavalid
		.custom_ip_bridge_s0_waitrequest                                  (mm_interconnect_0_custom_ip_bridge_s0_waitrequest),   //                                                           .waitrequest
		.custom_ip_bridge_s0_debugaccess                                  (mm_interconnect_0_custom_ip_bridge_s0_debugaccess),   //                                                           .debugaccess
		.onchip_memory2_0_s1_address                                      (mm_interconnect_0_onchip_memory2_0_s1_address),       //                                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                        (mm_interconnect_0_onchip_memory2_0_s1_write),         //                                                           .write
		.onchip_memory2_0_s1_readdata                                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),      //                                                           .readdata
		.onchip_memory2_0_s1_writedata                                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),     //                                                           .writedata
		.onchip_memory2_0_s1_byteenable                                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),    //                                                           .byteenable
		.onchip_memory2_0_s1_chipselect                                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),    //                                                           .chipselect
		.onchip_memory2_0_s1_clken                                        (mm_interconnect_0_onchip_memory2_0_s1_clken)          //                                                           .clken
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                    //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                  //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                   //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                  //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                 //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                  //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                 //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                  //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                 //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                 //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                     //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                   //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                   //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                   //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                  //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                  //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                     //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                   //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                  //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                  //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                    //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                  //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                   //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                  //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                 //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                  //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                 //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                  //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                 //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                 //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                     //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                   //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                   //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                   //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                  //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                  //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                         //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),              // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.lw_mm_bridge_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),              //                      lw_mm_bridge_reset_reset_bridge_in_reset.reset
		.lw_mm_bridge_s0_address                                             (mm_interconnect_1_lw_mm_bridge_s0_address),       //                                               lw_mm_bridge_s0.address
		.lw_mm_bridge_s0_write                                               (mm_interconnect_1_lw_mm_bridge_s0_write),         //                                                              .write
		.lw_mm_bridge_s0_read                                                (mm_interconnect_1_lw_mm_bridge_s0_read),          //                                                              .read
		.lw_mm_bridge_s0_readdata                                            (mm_interconnect_1_lw_mm_bridge_s0_readdata),      //                                                              .readdata
		.lw_mm_bridge_s0_writedata                                           (mm_interconnect_1_lw_mm_bridge_s0_writedata),     //                                                              .writedata
		.lw_mm_bridge_s0_burstcount                                          (mm_interconnect_1_lw_mm_bridge_s0_burstcount),    //                                                              .burstcount
		.lw_mm_bridge_s0_byteenable                                          (mm_interconnect_1_lw_mm_bridge_s0_byteenable),    //                                                              .byteenable
		.lw_mm_bridge_s0_readdatavalid                                       (mm_interconnect_1_lw_mm_bridge_s0_readdatavalid), //                                                              .readdatavalid
		.lw_mm_bridge_s0_waitrequest                                         (mm_interconnect_1_lw_mm_bridge_s0_waitrequest),   //                                                              .waitrequest
		.lw_mm_bridge_s0_debugaccess                                         (mm_interconnect_1_lw_mm_bridge_s0_debugaccess)    //                                                              .debugaccess
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                     (clk_clk),                                                             //                                  clk_0_clk.clk
		.custom_reset_synchronizer_clock_out_clk           (clk_hdmi_clk),                                                        //        custom_reset_synchronizer_clock_out.clk
		.hdmi_mm_bridge_reset_reset_bridge_in_reset_reset  (custom_reset_synchronizer_reset_out_reset),                           // hdmi_mm_bridge_reset_reset_bridge_in_reset.reset
		.lw_mm_bridge_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                                  //   lw_mm_bridge_reset_reset_bridge_in_reset.reset
		.lw_mm_bridge_m0_address                           (lw_mm_bridge_m0_address),                                             //                            lw_mm_bridge_m0.address
		.lw_mm_bridge_m0_waitrequest                       (lw_mm_bridge_m0_waitrequest),                                         //                                           .waitrequest
		.lw_mm_bridge_m0_burstcount                        (lw_mm_bridge_m0_burstcount),                                          //                                           .burstcount
		.lw_mm_bridge_m0_byteenable                        (lw_mm_bridge_m0_byteenable),                                          //                                           .byteenable
		.lw_mm_bridge_m0_read                              (lw_mm_bridge_m0_read),                                                //                                           .read
		.lw_mm_bridge_m0_readdata                          (lw_mm_bridge_m0_readdata),                                            //                                           .readdata
		.lw_mm_bridge_m0_readdatavalid                     (lw_mm_bridge_m0_readdatavalid),                                       //                                           .readdatavalid
		.lw_mm_bridge_m0_write                             (lw_mm_bridge_m0_write),                                               //                                           .write
		.lw_mm_bridge_m0_writedata                         (lw_mm_bridge_m0_writedata),                                           //                                           .writedata
		.lw_mm_bridge_m0_debugaccess                       (lw_mm_bridge_m0_debugaccess),                                         //                                           .debugaccess
		.arduino_gpio_s1_address                           (mm_interconnect_2_arduino_gpio_s1_address),                           //                            arduino_gpio_s1.address
		.arduino_gpio_s1_write                             (mm_interconnect_2_arduino_gpio_s1_write),                             //                                           .write
		.arduino_gpio_s1_readdata                          (mm_interconnect_2_arduino_gpio_s1_readdata),                          //                                           .readdata
		.arduino_gpio_s1_writedata                         (mm_interconnect_2_arduino_gpio_s1_writedata),                         //                                           .writedata
		.arduino_gpio_s1_chipselect                        (mm_interconnect_2_arduino_gpio_s1_chipselect),                        //                                           .chipselect
		.button_pio_s1_address                             (mm_interconnect_2_button_pio_s1_address),                             //                              button_pio_s1.address
		.button_pio_s1_write                               (mm_interconnect_2_button_pio_s1_write),                               //                                           .write
		.button_pio_s1_readdata                            (mm_interconnect_2_button_pio_s1_readdata),                            //                                           .readdata
		.button_pio_s1_writedata                           (mm_interconnect_2_button_pio_s1_writedata),                           //                                           .writedata
		.button_pio_s1_chipselect                          (mm_interconnect_2_button_pio_s1_chipselect),                          //                                           .chipselect
		.chip_id_read_mm_0_s0_read                         (mm_interconnect_2_chip_id_read_mm_0_s0_read),                         //                       chip_id_read_mm_0_s0.read
		.chip_id_read_mm_0_s0_readdata                     (mm_interconnect_2_chip_id_read_mm_0_s0_readdata),                     //                                           .readdata
		.cvo_reset_pio_s1_address                          (mm_interconnect_2_cvo_reset_pio_s1_address),                          //                           cvo_reset_pio_s1.address
		.cvo_reset_pio_s1_write                            (mm_interconnect_2_cvo_reset_pio_s1_write),                            //                                           .write
		.cvo_reset_pio_s1_readdata                         (mm_interconnect_2_cvo_reset_pio_s1_readdata),                         //                                           .readdata
		.cvo_reset_pio_s1_writedata                        (mm_interconnect_2_cvo_reset_pio_s1_writedata),                        //                                           .writedata
		.cvo_reset_pio_s1_chipselect                       (mm_interconnect_2_cvo_reset_pio_s1_chipselect),                       //                                           .chipselect
		.dipsw_pio_s1_address                              (mm_interconnect_2_dipsw_pio_s1_address),                              //                               dipsw_pio_s1.address
		.dipsw_pio_s1_write                                (mm_interconnect_2_dipsw_pio_s1_write),                                //                                           .write
		.dipsw_pio_s1_readdata                             (mm_interconnect_2_dipsw_pio_s1_readdata),                             //                                           .readdata
		.dipsw_pio_s1_writedata                            (mm_interconnect_2_dipsw_pio_s1_writedata),                            //                                           .writedata
		.dipsw_pio_s1_chipselect                           (mm_interconnect_2_dipsw_pio_s1_chipselect),                           //                                           .chipselect
		.gpio_0_a_s1_address                               (mm_interconnect_2_gpio_0_a_s1_address),                               //                                gpio_0_a_s1.address
		.gpio_0_a_s1_write                                 (mm_interconnect_2_gpio_0_a_s1_write),                                 //                                           .write
		.gpio_0_a_s1_readdata                              (mm_interconnect_2_gpio_0_a_s1_readdata),                              //                                           .readdata
		.gpio_0_a_s1_writedata                             (mm_interconnect_2_gpio_0_a_s1_writedata),                             //                                           .writedata
		.gpio_0_a_s1_chipselect                            (mm_interconnect_2_gpio_0_a_s1_chipselect),                            //                                           .chipselect
		.gpio_0_b_s1_address                               (mm_interconnect_2_gpio_0_b_s1_address),                               //                                gpio_0_b_s1.address
		.gpio_0_b_s1_write                                 (mm_interconnect_2_gpio_0_b_s1_write),                                 //                                           .write
		.gpio_0_b_s1_readdata                              (mm_interconnect_2_gpio_0_b_s1_readdata),                              //                                           .readdata
		.gpio_0_b_s1_writedata                             (mm_interconnect_2_gpio_0_b_s1_writedata),                             //                                           .writedata
		.gpio_0_b_s1_chipselect                            (mm_interconnect_2_gpio_0_b_s1_chipselect),                            //                                           .chipselect
		.gpio_1_a_s1_address                               (mm_interconnect_2_gpio_1_a_s1_address),                               //                                gpio_1_a_s1.address
		.gpio_1_a_s1_write                                 (mm_interconnect_2_gpio_1_a_s1_write),                                 //                                           .write
		.gpio_1_a_s1_readdata                              (mm_interconnect_2_gpio_1_a_s1_readdata),                              //                                           .readdata
		.gpio_1_a_s1_writedata                             (mm_interconnect_2_gpio_1_a_s1_writedata),                             //                                           .writedata
		.gpio_1_a_s1_chipselect                            (mm_interconnect_2_gpio_1_a_s1_chipselect),                            //                                           .chipselect
		.gpio_1_b_s1_address                               (mm_interconnect_2_gpio_1_b_s1_address),                               //                                gpio_1_b_s1.address
		.gpio_1_b_s1_write                                 (mm_interconnect_2_gpio_1_b_s1_write),                                 //                                           .write
		.gpio_1_b_s1_readdata                              (mm_interconnect_2_gpio_1_b_s1_readdata),                              //                                           .readdata
		.gpio_1_b_s1_writedata                             (mm_interconnect_2_gpio_1_b_s1_writedata),                             //                                           .writedata
		.gpio_1_b_s1_chipselect                            (mm_interconnect_2_gpio_1_b_s1_chipselect),                            //                                           .chipselect
		.hdmi_mm_bridge_s0_address                         (mm_interconnect_2_hdmi_mm_bridge_s0_address),                         //                          hdmi_mm_bridge_s0.address
		.hdmi_mm_bridge_s0_write                           (mm_interconnect_2_hdmi_mm_bridge_s0_write),                           //                                           .write
		.hdmi_mm_bridge_s0_read                            (mm_interconnect_2_hdmi_mm_bridge_s0_read),                            //                                           .read
		.hdmi_mm_bridge_s0_readdata                        (mm_interconnect_2_hdmi_mm_bridge_s0_readdata),                        //                                           .readdata
		.hdmi_mm_bridge_s0_writedata                       (mm_interconnect_2_hdmi_mm_bridge_s0_writedata),                       //                                           .writedata
		.hdmi_mm_bridge_s0_burstcount                      (mm_interconnect_2_hdmi_mm_bridge_s0_burstcount),                      //                                           .burstcount
		.hdmi_mm_bridge_s0_byteenable                      (mm_interconnect_2_hdmi_mm_bridge_s0_byteenable),                      //                                           .byteenable
		.hdmi_mm_bridge_s0_readdatavalid                   (mm_interconnect_2_hdmi_mm_bridge_s0_readdatavalid),                   //                                           .readdatavalid
		.hdmi_mm_bridge_s0_waitrequest                     (mm_interconnect_2_hdmi_mm_bridge_s0_waitrequest),                     //                                           .waitrequest
		.hdmi_mm_bridge_s0_debugaccess                     (mm_interconnect_2_hdmi_mm_bridge_s0_debugaccess),                     //                                           .debugaccess
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_2_jtag_uart_avalon_jtag_slave_address),               //                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_2_jtag_uart_avalon_jtag_slave_write),                 //                                           .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_2_jtag_uart_avalon_jtag_slave_read),                  //                                           .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_2_jtag_uart_avalon_jtag_slave_readdata),              //                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_2_jtag_uart_avalon_jtag_slave_writedata),             //                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_2_jtag_uart_avalon_jtag_slave_waitrequest),           //                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_2_jtag_uart_avalon_jtag_slave_chipselect),            //                                           .chipselect
		.led_pio_s1_address                                (mm_interconnect_2_led_pio_s1_address),                                //                                 led_pio_s1.address
		.led_pio_s1_write                                  (mm_interconnect_2_led_pio_s1_write),                                  //                                           .write
		.led_pio_s1_readdata                               (mm_interconnect_2_led_pio_s1_readdata),                               //                                           .readdata
		.led_pio_s1_writedata                              (mm_interconnect_2_led_pio_s1_writedata),                              //                                           .writedata
		.led_pio_s1_chipselect                             (mm_interconnect_2_led_pio_s1_chipselect),                             //                                           .chipselect
		.locked_pio_s1_address                             (mm_interconnect_2_locked_pio_s1_address),                             //                              locked_pio_s1.address
		.locked_pio_s1_readdata                            (mm_interconnect_2_locked_pio_s1_readdata),                            //                                           .readdata
		.pll_reset_pio_s1_address                          (mm_interconnect_2_pll_reset_pio_s1_address),                          //                           pll_reset_pio_s1.address
		.pll_reset_pio_s1_write                            (mm_interconnect_2_pll_reset_pio_s1_write),                            //                                           .write
		.pll_reset_pio_s1_readdata                         (mm_interconnect_2_pll_reset_pio_s1_readdata),                         //                                           .readdata
		.pll_reset_pio_s1_writedata                        (mm_interconnect_2_pll_reset_pio_s1_writedata),                        //                                           .writedata
		.pll_reset_pio_s1_chipselect                       (mm_interconnect_2_pll_reset_pio_s1_chipselect),                       //                                           .chipselect
		.pll_stream_reconfig_mgmt_avalon_slave_address     (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_address),     //      pll_stream_reconfig_mgmt_avalon_slave.address
		.pll_stream_reconfig_mgmt_avalon_slave_write       (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_write),       //                                           .write
		.pll_stream_reconfig_mgmt_avalon_slave_read        (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_read),        //                                           .read
		.pll_stream_reconfig_mgmt_avalon_slave_readdata    (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_readdata),    //                                           .readdata
		.pll_stream_reconfig_mgmt_avalon_slave_writedata   (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_writedata),   //                                           .writedata
		.pll_stream_reconfig_mgmt_avalon_slave_byteenable  (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_byteenable),  //                                           .byteenable
		.pll_stream_reconfig_mgmt_avalon_slave_waitrequest (mm_interconnect_2_pll_stream_reconfig_mgmt_avalon_slave_waitrequest), //                                           .waitrequest
		.sysid_qsys_control_slave_address                  (mm_interconnect_2_sysid_qsys_control_slave_address),                  //                   sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                 (mm_interconnect_2_sysid_qsys_control_slave_readdata)                  //                                           .readdata
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.custom_reset_synchronizer_clock_out_clk          (clk_hdmi_clk),                                                //        custom_reset_synchronizer_clock_out.clk
		.hdmi_mm_bridge_reset_reset_bridge_in_reset_reset (custom_reset_synchronizer_reset_out_reset),                   // hdmi_mm_bridge_reset_reset_bridge_in_reset.reset
		.hdmi_mm_bridge_m0_address                        (hdmi_mm_bridge_m0_address),                                   //                          hdmi_mm_bridge_m0.address
		.hdmi_mm_bridge_m0_waitrequest                    (hdmi_mm_bridge_m0_waitrequest),                               //                                           .waitrequest
		.hdmi_mm_bridge_m0_burstcount                     (hdmi_mm_bridge_m0_burstcount),                                //                                           .burstcount
		.hdmi_mm_bridge_m0_byteenable                     (hdmi_mm_bridge_m0_byteenable),                                //                                           .byteenable
		.hdmi_mm_bridge_m0_read                           (hdmi_mm_bridge_m0_read),                                      //                                           .read
		.hdmi_mm_bridge_m0_readdata                       (hdmi_mm_bridge_m0_readdata),                                  //                                           .readdata
		.hdmi_mm_bridge_m0_readdatavalid                  (hdmi_mm_bridge_m0_readdatavalid),                             //                                           .readdatavalid
		.hdmi_mm_bridge_m0_write                          (hdmi_mm_bridge_m0_write),                                     //                                           .write
		.hdmi_mm_bridge_m0_writedata                      (hdmi_mm_bridge_m0_writedata),                                 //                                           .writedata
		.hdmi_mm_bridge_m0_debugaccess                    (hdmi_mm_bridge_m0_debugaccess),                               //                                           .debugaccess
		.alt_vip_cl_cvo_hdmi_control_address              (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_address),       //                alt_vip_cl_cvo_hdmi_control.address
		.alt_vip_cl_cvo_hdmi_control_write                (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_write),         //                                           .write
		.alt_vip_cl_cvo_hdmi_control_read                 (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_read),          //                                           .read
		.alt_vip_cl_cvo_hdmi_control_readdata             (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_readdata),      //                                           .readdata
		.alt_vip_cl_cvo_hdmi_control_writedata            (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_writedata),     //                                           .writedata
		.alt_vip_cl_cvo_hdmi_control_byteenable           (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_byteenable),    //                                           .byteenable
		.alt_vip_cl_cvo_hdmi_control_readdatavalid        (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_readdatavalid), //                                           .readdatavalid
		.alt_vip_cl_cvo_hdmi_control_waitrequest          (mm_interconnect_3_alt_vip_cl_cvo_hdmi_control_waitrequest),   //                                           .waitrequest
		.alt_vip_cl_vfb_hdmi_control_address              (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_address),       //                alt_vip_cl_vfb_hdmi_control.address
		.alt_vip_cl_vfb_hdmi_control_write                (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_write),         //                                           .write
		.alt_vip_cl_vfb_hdmi_control_read                 (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_read),          //                                           .read
		.alt_vip_cl_vfb_hdmi_control_readdata             (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_readdata),      //                                           .readdata
		.alt_vip_cl_vfb_hdmi_control_writedata            (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_writedata),     //                                           .writedata
		.alt_vip_cl_vfb_hdmi_control_byteenable           (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_byteenable),    //                                           .byteenable
		.alt_vip_cl_vfb_hdmi_control_readdatavalid        (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_readdatavalid), //                                           .readdatavalid
		.alt_vip_cl_vfb_hdmi_control_waitrequest          (mm_interconnect_3_alt_vip_cl_vfb_hdmi_control_waitrequest)    //                                           .waitrequest
	);

	soc_system_mm_interconnect_4 mm_interconnect_4 (
		.clk_0_clk_clk                                      (clk_clk),                                              //                                    clk_0_clk.clk
		.custom_ip_bridge_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   // custom_ip_bridge_reset_reset_bridge_in_reset.reset
		.custom_ip_bridge_m0_address                        (custom_ip_bridge_m0_address),                          //                          custom_ip_bridge_m0.address
		.custom_ip_bridge_m0_waitrequest                    (custom_ip_bridge_m0_waitrequest),                      //                                             .waitrequest
		.custom_ip_bridge_m0_burstcount                     (custom_ip_bridge_m0_burstcount),                       //                                             .burstcount
		.custom_ip_bridge_m0_byteenable                     (custom_ip_bridge_m0_byteenable),                       //                                             .byteenable
		.custom_ip_bridge_m0_read                           (custom_ip_bridge_m0_read),                             //                                             .read
		.custom_ip_bridge_m0_readdata                       (custom_ip_bridge_m0_readdata),                         //                                             .readdata
		.custom_ip_bridge_m0_readdatavalid                  (custom_ip_bridge_m0_readdatavalid),                    //                                             .readdatavalid
		.custom_ip_bridge_m0_write                          (custom_ip_bridge_m0_write),                            //                                             .write
		.custom_ip_bridge_m0_writedata                      (custom_ip_bridge_m0_writedata),                        //                                             .writedata
		.custom_ip_bridge_m0_debugaccess                    (custom_ip_bridge_m0_debugaccess),                      //                                             .debugaccess
		.ctrl_register_s1_address                           (mm_interconnect_4_ctrl_register_s1_address),           //                             ctrl_register_s1.address
		.ctrl_register_s1_write                             (mm_interconnect_4_ctrl_register_s1_write),             //                                             .write
		.ctrl_register_s1_readdata                          (mm_interconnect_4_ctrl_register_s1_readdata),          //                                             .readdata
		.ctrl_register_s1_writedata                         (mm_interconnect_4_ctrl_register_s1_writedata),         //                                             .writedata
		.ctrl_register_s1_chipselect                        (mm_interconnect_4_ctrl_register_s1_chipselect),        //                                             .chipselect
		.lfsr_reset_value_reg_s1_address                    (mm_interconnect_4_lfsr_reset_value_reg_s1_address),    //                      lfsr_reset_value_reg_s1.address
		.lfsr_reset_value_reg_s1_write                      (mm_interconnect_4_lfsr_reset_value_reg_s1_write),      //                                             .write
		.lfsr_reset_value_reg_s1_readdata                   (mm_interconnect_4_lfsr_reset_value_reg_s1_readdata),   //                                             .readdata
		.lfsr_reset_value_reg_s1_writedata                  (mm_interconnect_4_lfsr_reset_value_reg_s1_writedata),  //                                             .writedata
		.lfsr_reset_value_reg_s1_chipselect                 (mm_interconnect_4_lfsr_reset_value_reg_s1_chipselect), //                                             .chipselect
		.random_s1_address                                  (mm_interconnect_4_random_s1_address),                  //                                    random_s1.address
		.random_s1_readdata                                 (mm_interconnect_4_random_s1_readdata)                  //                                             .readdata
	);

	soc_system_mm_interconnect_5 mm_interconnect_5 (
		.hps_0_h2f_user0_clock_clk                                          (hps_0_h2f_user0_clock_clk),                             //                                        hps_0_h2f_user0_clock.clk
		.alt_vip_cl_vfb_hdmi_mem_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                        //          alt_vip_cl_vfb_hdmi_mem_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                    // hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.alt_vip_cl_vfb_hdmi_mem_master_rd_address                          (alt_vip_cl_vfb_hdmi_mem_master_rd_address),             //                            alt_vip_cl_vfb_hdmi_mem_master_rd.address
		.alt_vip_cl_vfb_hdmi_mem_master_rd_waitrequest                      (alt_vip_cl_vfb_hdmi_mem_master_rd_waitrequest),         //                                                             .waitrequest
		.alt_vip_cl_vfb_hdmi_mem_master_rd_burstcount                       (alt_vip_cl_vfb_hdmi_mem_master_rd_burstcount),          //                                                             .burstcount
		.alt_vip_cl_vfb_hdmi_mem_master_rd_read                             (alt_vip_cl_vfb_hdmi_mem_master_rd_read),                //                                                             .read
		.alt_vip_cl_vfb_hdmi_mem_master_rd_readdata                         (alt_vip_cl_vfb_hdmi_mem_master_rd_readdata),            //                                                             .readdata
		.alt_vip_cl_vfb_hdmi_mem_master_rd_readdatavalid                    (alt_vip_cl_vfb_hdmi_mem_master_rd_readdatavalid),       //                                                             .readdatavalid
		.hps_0_f2h_sdram0_data_address                                      (mm_interconnect_5_hps_0_f2h_sdram0_data_address),       //                                        hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                        (mm_interconnect_5_hps_0_f2h_sdram0_data_write),         //                                                             .write
		.hps_0_f2h_sdram0_data_read                                         (mm_interconnect_5_hps_0_f2h_sdram0_data_read),          //                                                             .read
		.hps_0_f2h_sdram0_data_readdata                                     (mm_interconnect_5_hps_0_f2h_sdram0_data_readdata),      //                                                             .readdata
		.hps_0_f2h_sdram0_data_writedata                                    (mm_interconnect_5_hps_0_f2h_sdram0_data_writedata),     //                                                             .writedata
		.hps_0_f2h_sdram0_data_burstcount                                   (mm_interconnect_5_hps_0_f2h_sdram0_data_burstcount),    //                                                             .burstcount
		.hps_0_f2h_sdram0_data_byteenable                                   (mm_interconnect_5_hps_0_f2h_sdram0_data_byteenable),    //                                                             .byteenable
		.hps_0_f2h_sdram0_data_readdatavalid                                (mm_interconnect_5_hps_0_f2h_sdram0_data_readdatavalid), //                                                             .readdatavalid
		.hps_0_f2h_sdram0_data_waitrequest                                  (mm_interconnect_5_hps_0_f2h_sdram0_data_waitrequest)    //                                                             .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq), // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq), // receiver5.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (0),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (0),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (0),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk   (clk_clk),                            // in_clk_0.clk
		.in_rst_0_reset (rst_controller_001_reset_out_reset), // in_rst_0.reset
		.in_0_data      (altchip_id_0_output_data),           //     in_0.data
		.in_0_valid     (altchip_id_0_output_valid),          //         .valid
		.out_0_data     (avalon_st_adapter_out_0_data),       //    out_0.data
		.out_0_ready    (avalon_st_adapter_out_0_ready)       //         .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (custom_reset_synchronizer_reset_out_reset), // reset_in0.reset
		.clk            (hps_0_h2f_user0_clock_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),            // reset_out.reset
		.reset_req      (),                                          // (terminated)
		.reset_req_in0  (1'b0),                                      // (terminated)
		.reset_in1      (1'b0),                                      // (terminated)
		.reset_req_in1  (1'b0),                                      // (terminated)
		.reset_in2      (1'b0),                                      // (terminated)
		.reset_req_in2  (1'b0),                                      // (terminated)
		.reset_in3      (1'b0),                                      // (terminated)
		.reset_req_in3  (1'b0),                                      // (terminated)
		.reset_in4      (1'b0),                                      // (terminated)
		.reset_req_in4  (1'b0),                                      // (terminated)
		.reset_in5      (1'b0),                                      // (terminated)
		.reset_req_in5  (1'b0),                                      // (terminated)
		.reset_in6      (1'b0),                                      // (terminated)
		.reset_req_in6  (1'b0),                                      // (terminated)
		.reset_in7      (1'b0),                                      // (terminated)
		.reset_req_in7  (1'b0),                                      // (terminated)
		.reset_in8      (1'b0),                                      // (terminated)
		.reset_req_in8  (1'b0),                                      // (terminated)
		.reset_in9      (1'b0),                                      // (terminated)
		.reset_req_in9  (1'b0),                                      // (terminated)
		.reset_in10     (1'b0),                                      // (terminated)
		.reset_req_in10 (1'b0),                                      // (terminated)
		.reset_in11     (1'b0),                                      // (terminated)
		.reset_req_in11 (1'b0),                                      // (terminated)
		.reset_in12     (1'b0),                                      // (terminated)
		.reset_req_in12 (1'b0),                                      // (terminated)
		.reset_in13     (1'b0),                                      // (terminated)
		.reset_req_in13 (1'b0),                                      // (terminated)
		.reset_in14     (1'b0),                                      // (terminated)
		.reset_req_in14 (1'b0),                                      // (terminated)
		.reset_in15     (1'b0),                                      // (terminated)
		.reset_req_in15 (1'b0)                                       // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (rst_controller_002_reset_out_reset),     // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.reset_in1      (por_reset_reset),                    // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (rst_controller_002_reset_out_reset),       // reset_in0.reset
		.reset_in1      (cvo_reset_pio_external_connection_export), // reset_in1.reset
		.clk            (),                                         //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                         // (terminated)
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (hps_0_h2f_user1_clock_clk),          //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (hps_0_h2f_user0_clock_clk),          //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign hps_0_h2f_reset_reset_n = ~rst_controller_004_reset_out_reset;

endmodule
