��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P�:dG�!�y��8�՗T�{��9l�g�R1�:�9:{�#B�u�v�rG#\��k��u�P��IB4�փ<�:bS�2��T�%��������
ȕ?�P���$+����(�iό�et��&�]���|{4��A�I�e�A*C��6@����rGV:�w�xOK�P��+���Yï�ҏ`P(~��ާ�υ�Aa-zQ�t����� �6�k��U���nI��G�9�"�O��}ń�=+_nГ��!�3V.�>��kpn�o���7�	�?b.�\�bp����K�]�r^��������x%�� ���4��G�r����+T��|�!GR��p��E@�h��{��֙%�{�=����#��Q�������0�Wj��՗'�����=�*�N�o��ӝ��b��M-=����!vq�x�D1�B���5�ٳB�_,֧'6��v�F>y ��J�29��%�� g����yT� �d|�=/�S���s\O�5�|!�q7UC���9�Pה[��&���ƈ�W/���]?x�,�\p B��_'i��Hj�F.��C��]Ȣ�:��j�q�c8l���l1YI��>A4��a��A'>k�"l�6���<76�R����]ؼ�e��$�An�#��Z����x�3�f�����Q�
>�"�#2�C�U�ee��G��*[�JX�g�2�=/�Z��UEjȻ1�pE��B���(LA���j��NTr��I�c�t��`���)��}�R=�rT��u��\��C�7;��먥$�g2G�o�}����G?������NqO-��	5/^x�Ŝ�T�R��"_��� d�)��z�M`.�F ��:�x{I�v����w`����zsɕ3k����=w� *ܳ5�8�"]�:C�
Y�B�\�'��$&{j(- �l���f��<�jY;�.�A�Ʌ6N��)�]f���ϡ�Lob�A�+}BI��M��B7P�٠T~�k����~F(��3�e��L3Ū�Ⱦ�}j�n�Z�����8��?*�x��J
��E��v`,�Q�����㦑?b�ɳ�d�Zٹ�����PVL�̓M"�i���F�Έ����? �F�Pl4�:e��q,����C�m2�p]�?�8�D?��В[�Kx9HnI��Bs%jd��$qG�u��dBV&q��u �#�����b@%k��$���|+�2p�pC�8�bw=k?Hc[w.ǩ
#���q����f�{)Ad��!��vw�-���H�E�#�6�B����kU�P:*�L���C��a$�w���7a�◼�b��"�n�9�vu��A> ���y淘}��}� �F�@W||��ȓ�Ӝ1�.$�$��᯽1m�����ѽ��r6�f�$p7�`g���@�|����|��o�TJ�۲#�IڧM\g*��k���}mB��&:�*��V�l%ks�:<��L=3�?�Q�� ��7w}�,�F�{*���]��&����~��<�>��/F���9Z�(�>�{�n�v�A׸w���q�m���b���+|3j*J���3Ǯ��bu���/s��I�Y$،ktw�<��ބO YSV�H1&���.2:�!��m�z/X	�3�R�>1q�}�<v�L���DD�elސ�I\����;;Y�\�D��)�G�jC*;*��-=�g�$
mBm`d;9����ϝ�⎴�H�鷈_��� ���2�q�@.�]��H���~���tm�À�3[�*)��N�lK�p�us�=���!���fP���gdsTn�a�.{��Yr`^���)t˗�e���B\¡��F|�7yi>N��K�԰�"9����2 ��h$�~gU���
�7<�L�Y����+�t��V��兡.�����yt�������2��d���K0�+�S�J6X��Qi�B� <��J�t�O��ٱ1N�Cp�_\؟��[���g�b�R�x�����2�L@��Tut ��Mۼ���N�k}�}������^������>p�9���8�m#����"�z��DQZdG��RVb�]8����Ǖ/P��� �?�?H*�ɪ���ţ�IV��n�?�6=Y)H�c�4u7�	� /�8��W7���Ww��؜Y���A�R�Et�?����Ni����$U]��^�a0Gؗ��I�Դ0��0MY�7������s%N���u�c���냚�7����b�b7&��Ф�N�8���e��RČOn/���T��G�dc��}�'��-iG;��O7�Ͱ�a�_��B��y0a��F[(/i�q�&me�\r�J���O��?���Z�ߌ?�;C�40��|M�����RP#�8�&)p���۱ڡ*ȍ�����1i�Y�o�j$y"B��h���_Ƶ������U��M_�ҫ`Z��&����a$��"�a�����g���W�d, �L)}FH� nڜ󐓢Z��0��00�tnJ-{$�j�#�3��%h�J�/� qc6ތy:w����C
[㞲�+�9�j�バ �y@Wr�<w�d��O�t&�)�������jBх��/����U\a�+$AE)GM�����X(��C6yO���Ę�x������J�;NIC���|��L����LD�[�����n�g�45Oǂ`��dY0��?4#��`ŝ ��nm7P4Ɩ����9��ī�on�*ox�ܜ��]e�x���D�b�qO�e�B�'�E"D뒳���ЈC�悈��m@܇��B�/̉�L��!�&jR)��9NZ�G!�t���#��I����&�=���+������G�c߶��p��f��/R��p�W^�QfJF^+�7j����#,ߕ3R�܈��[l�>Z�Y���M�4ٚ���Sa�%���n����c�N��9�#�а��D��D}�z����yw<��&c��4�z�I�w��5(��Iz���-ęҖ�o�?=�/�� cJ�+?�!����*�S<^`���4�qV�,�����}n�Kч���Z���;����0�����qN��Vdz���E���/Fm?���\#��<[2�DA��B�Jߦ�����{"�B���4�R��`������v��3�^�7���kIa�=v�ϓ��4���#0Oأ��t2|�EJ�����D|���d%V-xp�����K�r.��x���F�[=�g��dh�@.���/Hu�P�?�s�GL>��\�~��[��q`?�r�k0yB���oR�/&�o2�)��s���7�[_��2�URb���4/���5>��Ch8�2|�v���[��;3Gؼ��=w���� f�sɜ�0���$�x �����fњq.��c�"ֺҨ=�
�l�^��o����g�ٸ��R,��!!l7 c5�	�]����RD-~��M��b��}�D����������y' ��ٳ�S
�B�L7R^��f~1�D]����.�,��C�"O�,m2�ƖP���&�4����c� ��đ}Q8���z���A�+ݽK�������M�[(۬�ȸ�PaC��0��<��wq�+uX�� ��AM��@��L^92�<N�Fɂ3Q�}5py= �nȸ��v�F뀼�����D�܋�X�яa� �d��E�d_,�8Օ�K�[��u��6�$�S���[����<Z�\��Ĩ�?��Yo)�P=��I{�ӟ
c�֢�%��+10�|M��g%�w���Լ$!��sG����A�y�n/te�Eu� @��×05���j���eQR�tr��z�E�`��O�g���1�ߤ3���5�oki���n7ay4�S�Q竨�Ԙ޺�S9\^Z���o���7�Yro��w��c����(LZ2���R����1#51�0dqe�nGvՔQx�&�)���T�[�h�:<�I�a�Q��Qb��=�T�pft�0t�ΊL��ڹp��^%W�mƴL� \�e�Y�Cy�-?D����c��ʊ�:�sXZ�|v�%�v��/��7-2}f���ؐ2\ �|
�}<wњ0�7ܠ���b,�oM}���6��sz�eIi�v���,~T�ɨx��c��Ϩ�_-Z����t�&r��JA��j}#�Y���w�AIf�B>��*� �L�F�Ҽ��)�v��r��ON(��*��*tp��],�i�{���b��| �����:{Wl��-��<��Ï<��i�98
�Hjg5L�표��Z���]�[[��eޠ��L։��Y��;��:毖������9ǷϵvǷJ~L4a���͓B���6��@ٲ㼅oȄ��(Q��"���p�Gk��I�lH�"&���!L�
�}9"��q%;���8�ށ�h�*�l<q��X6jDn�3��	,j��S�2U�=R�-�!�y!���[hx\��S�������i��pk��X���$K
�֩rۥF��o�p���C����3s��	*fzhם�W��Τ'����0?�cd@��e��/��5[>q�8�a�|�%��}$��9Z��wl��Ь;�z�XΫ�y����8f;��d�W�6� �+vL���Z%�������J�QũT�"��)'��s�x���Bpyu��e�Cg��#\))��V�;g��<�k2E��Bg��Ŵ$�^�e �#��T"��'U��1�<�Z9K�����"-{���q�\������W��H-՞(��j�ic[� f]�5N�\!25��X��_8��� �3�;�07U�1�Y@=������2���C��}��&f-�,��u\�0��	�p�4oI��E�^:}��v���V�����[\�8�е	l��%�q��KpWO���&��zCۇW�3��gq1��n����V�-"g��քMNa��OhO��F�z�������"j)���h(��W�"�@`�85�,��,����Fx����U�\0�W�7���ܓE»mnZF���͠��<
��g��LT�[q����t
{�E^9P\�'�B�0A�µq-�sȑ�DDb)�Al�����wuq7ce�7��o�5��.=���u�e��Lg��K�^pxմݭ�iz����V�����ͧ��P��_�B�z�����p~-��ɲlM�n�;	����	��P4�T;��do�
���|C��^<C�L�R6��"TOI�w���AL/�$ùB\�_%]��Ʋm[?8�fC��r��ΑIb��U����;x��*�]�����֏�p���֚�i�>��Y�+6�7`�6!�29��k}�#�)(�hcf �j��u���K���m`�x�Hy��X��C��ּ�D�˞��7j�q�<a��� 9�$��Y��yvc�d<�8��q,�$��"D�.8�+<G&�6xX9���%�����Q���(u���8h����3�TcX�1��
lӏ,��(YO�Qe	�S�ݛ�(���9}����`z�^�@psw� ȴ]�{��n�.ⷜWES*/��.pAc����)�q<�SS�c���A�|KE���� �t+޸��u(sxq��&s|؃���������u�u`����_���ЃV7��c�˴
@\�R=̄��=|�	TݳX�����ooB��/C�dq��^>m�������y��h��YH�G�{��B�K߾�ԕ3K�ݥ�����S�d+�c>��%��c�e�5F�������� Z�����W��~�0��t�`�!}.k�I�'���oA�Hc+\?�W
��3}��A�=�l����FA��$�C��g�7�^���bA���PU�ꗴyLM�yڒ�q7�0f�^o=zш���Y�]��+�4�u_���Fj�,���GX�Î	ʭJ_|�ӊ�jQT7qW��	p�7 �!:��GM�Aڎ-��L���g�7�gi�>��Z{�=k�f�_L GCOL��s��8����
icbχ�y9��MT��r�gm����k]r��4(�o��%��I���+~I�3SޕB�7���c?�$����P���4գ�{��#�׽�N@���[	����@�����ܟG���8B�=m8��g�@�=3�.��:�:�N��|�] �[�:��s�IW:���4H����(v���McƱ���{�^���O�?ImZ%]�rU6���Kz^�>��C%�aw�.����{�@��-1��8���0{Cm�Jˇ�3H&������)��#��ڐ�V ucl@����f)h�Q��2������%()��:*�b�#�v�G-p(��C��w}���h�w��tl��T�d�����Z��9V�Wo���)�@��Lrd��Z1�v��ܑ�!Ș�w���I��׃V���O�L�yW���F��FI	�$C��(���l��;�1]k��T5�1�%�������Pq��&ߩP����븂:�iJ��*&�	0s�cH��ɲfc�닽�y)�VHK�,L˓��dĭ� �j-@ָ����Ů6 �1&zxU3n��b9%-ÞM�R6�ed��������I^9l��V�g����b�7Q&������k�K	�wOf@��uogr�1���v|x�� ꓝ	�ޅ���`�=2 v(6�W����민�ב8K8g��V&����~L3y/���%Ӕ��^���8t��AF��-�8��˄��Æ@�Bo�b���{��.���ݔ����v�^�'�X��+�>�,�$��`$��L��f�4��}�˅���T�D�|���K�S_���[�k�bc�+8���	Lu��"��}���l �&T\��_(8E{��C�:�o�@��Q�JO���~)rz�=�nLmt���a��\��.�|�����~<��MT*�r2�´��7cn�R�0�%�/ԟ��rW�F`V���T���O1���gT�8�I�~S� '��MS��4�w:���N��3/�Yd�fQ}Z� �h��	'������ia�b��5����}3�!�Zk�;�+�m�\�L�%����|8P��-�c�G�Y��&	~�I���*"�N��GI/(��XQa���[�*@��c��Sc��-��y��~� ]�e�4������J����v`�q�h��\� ����>_x�B�^#[��彼t��o����ݙ�_���(�
�:��g�?���G�m?�1]�;:_��qR����P�\��H0�06ǚ:���+��n��ٳj40�ΝSg��[�b%�.�%�V��iO��t!?n���%X�N��i��־u�b{v66⊌ب��DA�Ş4ν�~ꨮ(Y�6y�9���jac:��w�1����"f̓k�"��fd��V4�+�V��*��Ҝ�J
�!�Wm^q�}y4{p�����V}��0-����q�&���劥䯏�7hT�H�ٚ��)Yv3�!ὃ�.,�`��.!�̕�A���9�lo������b@�\2��~M�N���_~o;�J�Q~�+�x��4RM�7��Rid`�
���|��Ҩ���w�)��!yƠ�*�������{���j��ok�w�Wg (�m��� �ݐ�l����T�M6ŒZ���4��l폐\s��t�`�\�/��Q��.y��[� ��(�8�|%˱8��䭥'��c�D롙W��t��ZL�G����9U�LgK��j��T����t�5�~uˤ��c3�V���F����:z�!��~�-�i9���ZUMlaT�������Q���c'�L�Ot�����%�}'=��Ҁx��|�6JWWI,~��s�ƫ,�˓B��j�:���ic O�}�湪ݣ�xoX��E#�ȹ֚�ZI7s��+7M��F���1IG����G1P��OQ���涪[G�o�~!ʫ܋m�L��훝h���	�#ܶ�19_�:΄U[��_�"Zl��ԯ*�GG�S�
�3��������>Xݡ\sZ8��Ue�f�l6��&>�r���5
__��6~�>׿7S��l���oa,+q�Q��v�FSJ������x��/'���g�k9��ې����8)7�g�٭Q=�SmM��DUñ���9��~L��aƏR����8U��3�6��T�����C���VL�@�LH��	�*<"�}��mhn};�^zՐ��Z*i������Fը?��E��Oo�@^~�ݕ3�It���n���7��6�.$7b��׼"jcoQ���?�A�Ẅ�w�jB-{����Pժ�(p��b&>R��<�s�W�J^�/�:����	BJ�p��	g6�3��*�
�\���,Ȧ�;J���`��Z+cB�(� Sy:|�~�؉E{������9�@��?��t���!Gj7v�O)��-�����L���JV<�3��/�0c@�W�ķ�L�c�r*�ٓ+��ѣ��'�Wu�j�f1�	�MOF����@���@����F�ܾN���q]�5)�i�v>Eh�)�p��q�����W�e��R1S� t���S�O���������u;������Tu����KiZ��<�-y�B�S�VO5�y�	�I*�sqbgx��}sK�8t��E)�;�>�7ŝA���Ԗ�s�.�\��e�$VF&��_-���d:�43�;�SW[R�/)ں
`��N]��{����ʈს��*�N���̃.s_V-��%�D�$��E	�ܴ��Dj�P�`���sӧ[i����6z����� D) iP�RȖLs1�?�1�:X65�����',h�.���؁���U�A���_K"�"{`F&����w�B�HP!D�.])b�֝����J�k��jp�f;���j�� �J��^����~�����^Z�0�u�B@�0YW����*�|٣�ڪ��r�ܜ�YQ�QN����v~��󚏽]1�~:��jB>k��G�R���`C����K��#����x��.%D���/T��^����Ų �nH��&u�Ez���[[�㫇��F�P�F�n�3 :V��ć�N�i���g!�J�bM��C2-�Z�œ� �vV9r,��rǧF�oV���>��a�ca��q���׵5���nDD��	�h����<����x�7E���. g����6"�w�:�|��Z�Qg�y���h���NF�w�c�=v��ģ��F��co�\h|W�Aд�*�A`*(��q;��H�Z]��B�hEs���\��('�+��O0�GЂ�G_���ѳ�):BxY���ô���Y��zLS8 �2�38�����ā=]d��P����t���)0�v�R1]a�1toqf�y�����Jȴq�KP'<�o������(pc�_�IW��X�HHЬ�9�*/8�� n�di����?ͼ¿�9�S�
)K����R>��J���~M��Ǆ�GN�`!
�mçI�wtCo�]�B,?ީÀ5:M��ǾbCl	5\��mv3�������h��u��k����%�@U���X�_�돵n-&މ��E���m�}6s��$�'�倻�/�K��DL�p�g&�m%�}T'��Q��{��k�H�b�+>C�-�!��I�5�Z޳���y�$B+�W�&�O���蟬=-"VE�@�ut��Y?э�qVn������s<�<;�� .R��A�����5��nJ"_m���<����7(2��s��}S��g4,����%��T!vm�P�����'�`C�x)�۳�k&�[V�����6Z��(Z	�����x�;W�8���gB� n���
}"v0L��')�`T7�}���,�:����{��<O�»�G�{��C�0���>hdV�Y�j�x��"��2�����	�5�TF�� �Լ'p�߆��j�Rӓ�.Ms����/#g�\7�K�w����+F�EP�.�Q�f&}�aI+��q�nq�O%_D�v[x�S�i���_$1�OP�0��:��zyj1��H?���JG��e\,Q/'�P��������E	�B�+��jR5���������&D�F��bE�f��N���}4���,q���}S��������}	����3�*��kv}������>-@a?=�q����<�<K��X5������Jj�?z ]������j�\�ޭ�(��p,��
{����oB�����c��{f�+S��3Lg��c��>���f�-I��}��ҍ�3�؈��.j{��f��f,i|5�/��j���놿,���V���6_@1NV��*��M05��-t��.���[����pO��3o���^�.��{�eH�#���n��՞�Tl!�pd�^4���NRD�$b�1���5C�a����L�ڕ���t����)EoTU]��-�����<'���]��e����+XpW������|_����y���B���\bj�դ��G|N#o=?I׿�;#��4eap��~�U���z�}܇oƱ6�A2_n6	��\���n| ���V��y˘��f{��2�ݕ��Ŗ��1���֯�bTn�1�u9�g߭����p��G������a���[��D�3R���}��7G��舛����6m��i"e5a��u�:�RVf�C��;��B^�U�)3�a�7j��d@u.5�f�;5��Y�"����26ሐ�7"�fl��+d>U!�Bs��L���F��W���]��r��~������ti��sC�s'׬�a4�)&�R-@�d8Ը�O�L������j���Yw��i��3�|�h�-pL�����_��
	拮�6{��N�:�H6��qȡ"Ѣ�I~���[̂V�)�(���U'����9
4R�{8���dҪ"o�`��!R�1�Cp�u�Z�
ZTs4��F>��b2��1)��Y��<���	��%���ƥ��9go��-�g���檓�p��jL��O����݁�
�h��Yn`���p��揧u�qY���􅬈���-ς�����E7��0x�?��:P�D�+!^� g)ɓ�`�<��NnXz1^��zB��`�ޏ����V={�M�҆x����t�ְ���v�6��6b�[�#X���%�$=�fN��Ѵ������nC�s��β���� =��;�Ԡ���}��I���"E�Q5k���RQ^�w�^�����u�{c:����.�v�8,�F��Q����zT�å�)��������ѼX,#�vgn�ߜ����$�뤰�{Wz�o9�x�'�S+=}n���SS1<$�1��������R/���ZXT�eA:>�}m"����N4�RA4����֩6�(��Vb"�m�G���ir�:R~}ӭ��XM��0��y�_�L-3�p!�N`�lT P=�	��'����y^��D�[��t��{)?��r��0h��Y��'ϛ�i$�Au������+S;��Z������C˦�R���ݶ�\j�3����$Qi�+����Re+��?x�dM��Lh)�d�5:����+�(���������04��&E l�.�QV ��<����+��(/Db�)R� ���+����<Gp1RKb�����4��\��
��~�����$:|�>���@W����s鐿V�����-��1?X�Da'��()����&����\z'ï ���6�r��_\��ت:Ӑi#�L�*���b��>+)D��	b�xW
����;B�B��ՊS5��!-����W!O������W��N��n�,\j���J�9g���^R
����g�c�mB[�B�s��b�AtK�G�ot#�\c��nA���`�ԸG������e�8��oG�ߜ@N���Lje�=>ꃪ/��)ԘzP���MU����vw퉎���E)Ugņ�5�(6�ޗ��AX!N)�=�w��.����d�r��SK��M��<��0N$�ِ��b��A�$Nr����}�6=�h�Ԫ9VO�uiMT�uL��t(�I��H�z�>׌{�'�>��*�ul���DtѿϮ��������w��ژ�C�1e-8����]�����S� ����S��࿒��*�T`ʹ�ZL���^�v$����vj��]~Z���)~c��Y����%�p1��M�͈׎N�f3ԟ�2*�w2�K��6`�Q�H��ޓ�B�B�<�N=��V�&�viF�G��d�?��!�.���\4�y��9�OL�"L8���S��M������,�h�z�6g��7p���΄�<�>�cE6d5�i��u�۸Yi+%��ǵ���("f�mo�1@"W��T��/G.��(����1�.�c�4Ϫ���K� Y�O]y�U� �R��󂷇Yf�����|Ih�Nf�/4����ǳ.)�F��ac��z��Bם�i�D�Q���t�z�Ƶ=Z%�ī���¢�T@L�#���������s�Yя��b7��g|�2��o�;�/����j�@�ϻI�<Z'O8^7.#�qY�IA����x�.�W�jU�1+�lv������'��[���|��p_NŎ��(���O,w�vб �]�F���%�yù�y�}~���3G�e\4W�_���Fe�ҩ؟��fJ](t#E6�#L�����;���oioΙ������NN���}J�/L*m
�LP(܍0b�X��ւK(����N>�p 8^x	��>���t9�b}M>7[L�Ex�Y>L�J�`H%�L<r����0��H�>ݪ��M�y37�oa��u-�
�Qӈ�ϸY}t�n.�%:{	��1g����j�.�T�ĪN'����;��(l�����D)�%%؋.��{ٷ�w_3��Ѫ�"�ƫM�Xf�����Lx�q*�Dg�EKɸ��Z\��G� >��l�����z?u��&��Ϳ��\AH{}dM� �ߣ6?��NMC�`�r�7�Y��8v��W�e*{�[׭{b�솂�����r������hͥ�����������@#��D�z�ۦ�*��`�1f�N>b#��4t�c�����{7�j�^���g��SD�Q�XH�A`�H�6�� ����GFIZ���?�,'��n��J�RԞfݎ>�M�Pl
��x=�������|� �_�����hS)�I G� ,�[�c� ���cD��M�\��D�"}���VI�ap��{�;�.�Zy��l���8=@-u'���{�n��z�ɽҗ-@�_8vȾ(�p��>�`���t�X�U�C������;�% �Z~�g�L;����D�.��59�!ś��CL3���y�<5w+�3S���l!�����o�NQHPVI&��׈�2�}(&�F1l�r�t�%���2����sk�o�T������nUʹ�_�y	���O�t���>H���/Қ#�]�E����5(m<��V|�b�'��ΐټ��O�+��@�:��J�"m���41p�*�z��ג�IG��A��l��M0�U����o��L���[�� |O�T�{�.�����=hgt��D�1���W� ��ވ*����I���A��F�Og=B��^H����׮S2��:gCC��P�Bh ���q��y��+�gK���־�a�+؀,3YE$���r=`k���
�i-�YȞȧ,�̹��2�ǎ��-�TJo���3�>��e����o���A�s-э�Mu|�E�Rd�,���H�T�D(_]���;���k�DY5��ϖaI��FL�� %a�ޞ��#�M�U\]brٱJՊK@��>Ώe������d}ūmu�	�1e��tS�ޡ�b���f�G�G�j6/k�`��4���?;^!�����e�{:��O�^���#�8wW�w��r��GqW�sI>�V���\�s��L!�0�-6~�ƖJ��R���%�'TY��W��ˉ����SAݹW�Qtd��l�!m�D k�Wͮ���O0t!���w?̈��V/�0(b-��N�?}a2�j����uHa)����s5�:�.��Ǎ�E,|����#}����`�[ќQ"ԍ�����&�	k��ŕ� �w0�f�'�|�$�G'����$;��� ��!��Y��Z ��5����:TAz���Y������,_<y�[0H�����4W}VA˚��i�e�������N�~/Z$s�����)�Y6uM����#�W�WY/)�aV��.ɇp���z�L�ʷ��.SD���%�6�%�5椮>+_b$���ob��Kg�.�k.:�U��e�
@��Q�z!a�	V�:���X�!Uk������1A�y��Al�-:x��4�`F�cER�J�9+�������ꜭW�Fg�<�]��@�|�@D�~�Џު�Ӌv#�����m��wi���>=�p�Ú�S<@�W�;bX'�(��fn�h��[�{��-AR���O��Q��{NC�x�O�M6#=/�J�"d���w
׹��t��p=�*.$}���?��T��ٴ�0�������!�y%
�C`3R�b�^�*��:�����r��E�,%�v����;�L#BO�WY����o#Lx� �,��{WT3i�5e�}{�W��;�%f���҈,Γ��J������M�O5��%�8��((YxH67+Խ�>r�Bk�\����3H����h�1�Ĺ2m �ef���W��U�G*<��C�u�P�+���{@ʱ������ѫ��Ĺâ�΢��,���x<�nty�	�� T��T��yT6��w��%�ړR��j����$.�Z$�c�v��Yk�I������8��X����2�=S��	�T}�}b�%������ҩX�
%!�1p��X�٧J��f�Ah�WI�^f9��Q"]c���l�7�\�=�k���'�b3S�<�����(�ni���UU⣩1�}|� �ƥ���!�L�8:*"%�l~�EC�^�Q�FB�ݭ��@��� Y6[a�_ ��H��_R����α{�IR�~v~���"1%%u���hmc�Wqy%6��R�+Ƌ㆓ȭZul<�����;d)��u�?�J"�g�(������6�d��׾`.4j�����A_�-K�|=���l&�G(_��sI����3t��"����Q#�M�Z2�z^���CB�w�FI�%<9<����A�A{�Xf�S�q%zC0��*�wxfwTQf��9փ����&�C�u��m��Xa|�� HKH3j�e��ۘ.X��D�W�D����b�|��Ƀ$��G�����P�
�a�u��%Z'��j����+O��ؤ8�o�7�Bu�o��G�y'a�Z9��r��6+�d2@gx��y��dL�U�M��;R6�|����v6�,���s�i��dM+	}���G������\g��+32`)1�A�Մ! ���l�W�]^�pTY�V��G�ՠU:4r���>Z�����I`opH�z.)�� �c9FO�򕻔w���L�u���1�́���������<4w��wv�"V�.4��X�T׭�,����l�r�Hch����bt`0������3!���6�3A�g���	�
�.�g0A%g$�����T���	]S!�{���{�s(�G�X���N�e��n�܅�Y�wh��;P�^4^j�>e�	��11�q���*����2{��<>�9� iF��D�\�a�+�6������]��{���kT�g2$���F�ٗ��>
$���i6�̕��|�n��ƣB��
�I��
,Ȯ�.&>X�<3�[������ʖ�i�L]�׍���k�R~�?��
�T������#bG��f9�g6��鲯E�U1�`���4�6]������jֹ�X�=���i���!�x`w��a^)n$��H5�͝{�+}���$����)�� �;��?]p�s�\���v�j6������!��9S��,�b�]!X���+X���:Ϲ�R)����Q#������~�\/�i��Ԍ'�W�q7i~]jV����3�l�3���)�7��w�`�׳Kw$	%U��k瀾�7Pfn��}Fy�獩$�!��gũ�_�~��'���V�~��j18!��[���[�G�W�?0�G���/��Ms��.g���KE@l�G���P�'��V�a��1�dU`!$�cޞ�@n�#F!����+��3ďL��S8҃�!=�?q��������iy�[\C��6��\�I!}�~��5�S���k	]P��*��8 %���Uyz� Ɋ�m�r>��E�=,��H�GÐb�dSZ~�V}2�a�N�&X�<skH�L���:&P��V؍"��!��P�/���|P�liH��"ZnHZ����"EQ���o��w�w��-X�`9z�]�Ƃ�]6.�:=c,�0�$��3��R��K��I�0Nz��{s*���kV͡,���<��f�O�+��7i
#�ĶWx��9[G!x8j�O" ,W�%�*:�A�~м��wό���܌.��[� ʇJ��q�))�vm���e�t��|'�Nk�ԉ�%�ҝ;ݼ�e��*a։:I��6�[�L8�k�UT�wx^�V�YB���Tƹ)����H@��W�O!��3��Ykm�&ݾs�o���{h�,wҳ1����M/� ����I�ľL�X��a�k�?}^~������u�*��=��?�t@v&��D�0!�v��=aN�z���γaßpۚ�dz���0�X��ͅ��vŻ�n�i�5h��Jn�u��F�N>�X��H�%E��ͺ�%�j7�u�� ��*P���v�<F*m�3�-�v�_K{����o��<aXH�i�-Ǒ'�h<]*��`�P;ѓJn�Դ'���rr�4�=��c������qќ:��lh�BV��u��2��|�tMl5$���3`��a��g�|�J&n�'�R��ʙ�K�4-��C��<�Z��5��5�kpq%�	���&�P���Ng`�fy��%uX��~h��b
>^`���|4Ĭ�3q\Iҝww�1G��,M����V8�]E�J-�y{/w�fs
�M���S^�(Yy�;���%��[�.Y��h(� �t`�;ϩ�(]��+ֹ2����t5iP檘���Ȗt@�x7l/�����ϲ��Xr�P7Gy� �v�<@�������iV!���u%_��fwIE�v�=� ��x"��.JUܲa{���z�V�Z��ұVV�a�h�)�N5
B�3�ɵ�]�_����s� �P����{�R����Y\M��E�!��F'/��,�E�� >�_�;�K'��v�Y	���g:���r�xip\���'���Y�b���K��u�Bt��<�F7��6*����K���W��Px�b8�����&�2�$r\y�v%%-B;B��Y4��9O!��e���P��|[�贯ƂP��-'/gƘ�nm�qJvDo!���4,R��3���k6ө�wJ�ƛ�"�s;��J*[=�푉
l[C�^h�r���&̑�P�����Lޟ�1�QHX��r��Ҙ4¤D�`$З������SR���8M9쑣����\�6Ř��C^�2��e�n~7��7�"A�w�ʪhz �=_���eX]嗧wp��U�#�VЖ����G@���"q�Y'\]�����R�B)?���Ɣ�%)�Y��U��w~'���k���B!1�U:�˂P`�i�J<Q<�S*��@�y�GxoN���	<M{���}hל��r�ˮ�(��%9�N�@>s^���̈Ȏ��e�7k������<���h?T�[�ɓ�h��h�e�r�`��I�"�ݿ�� V�\@]Zɔ�אg�Y̱o��g�5[M��#�vZ��n1�ڼ�Mcj�|��L��W8?��ڏ���%��jE�Y�� eu��2�[�۲�\e�*����ޚp1��[��9n~鳾�(�JS�0���!\�z�1Q���p��;�D�h�M�W�k$���o�� ;�ݦs��{�Nn욽�p��� ��K3ѧ�򖵣Q/
{�&ȏ@c�(m�5`9<�CO���F��qf��}C�~�p����/�C# �T�(R�8�lM%���*�@�ԾL���,�/�}��(�V:��/w�{��gN��H��p�T�h�jAO׎v~P��Sͮ~V��$�X���J806�H�(�7� ؉��p8�$�"����-�u�zז�/x;{���������(��_����$ː�4�NJ"
f ��6}�6^tdJItr�[��E� ڒ|���Ez�D���m���yм�N `A9:>0e,�?���Jck�����nv$�c������?���p������#`��`�����������b��D'��bG�jf|k ����э߸�E%��?���
����4�>m�F���*^������}i¾	��$r8�����+s;o�:e	2�W�ڄ!�nt��8��0i��xwT�y��G��"'������_TJ���6��;/]5�?�tt���G=%HNeC Lp G���e;?���
5��؋�=u�iڠ�!4�-U~�?⚬E�{����?ӌw��c(蜱�@�fjd�=����� |}`����j���B=���P�=�6��uپ5�1ᯒ�G�=>x�I�H(rﰊЉ��g����X/�V�l�B��<��!(�G?��#ڵ	ÓiV)�@�x`�o݀��u�(1$ŭ���L���b���T8j@�p�"L-��Flx���Ⳇ�f��A]�Q�Ru**]��ܰ�|xG,pfh�'�U;sR�U�b�|��;�cv����#J��~�i~��2�T-ϵua��O�)���>�_������ӻ*��S �B�z�i��h���Pi���������5+��,Iۯ�wg�?Ҕ��ա|�L�w�_��6K��I - !%�Y$MjD�X�J�<"���k�<99��/R��
"ŏ�Gżn���vB����(Lݽ#�nu9��D���ߦ�t�r�s���]�>D/.N�����,���b����d��e�M�b��up���5P�&�Kǝ/�g1Js,������h�$e c���;l�TM��G���a�i�<��9x��GM_�y+z;�����H�4����|��.�-ӟ(���"��&�rH�Ms��׉G����*{�d���U:��{��F)Y�M���T2� I�<$Ri9)�a���4B�������┾`8Gc¾�岚�
����=�5.���\��k-}X��F���4H��B+'cc�|�������U�+��	���5�NByȍN���.�[�ji����+���'D�����e�$_`A8t��k���s~�S,X��Q�z]�A�����O���0<�3%�`51>�p�
�s��3����rl�Z��m;��'���$ql|"����	���/��p�b��Tɡ�l�G��p����O� �^8d�E�f7YJn���q�C�d3L�Py���)����=Z������^۴���H�DO��qb�S�Ka9IELD����6����^D�G`�!	�G��	�W}Bݦs����y��B4�,���	��<��C��ON�Uy�����?���rF�0����f��}��d�o��7T����Y!���&b^K�����V {� �*w�on?2����\Y�n�$`~��8�[��	ͬ�����7��8E4�l�&���{B��3�4F)|ā�'��y*��������r#���f�fl=�x:��F�Ź��ٷ�KX}���w��O)��%b�����.��=ٯ��R66�&�ƗI�HT�J�1F���cesZ����\�����;(RH^K{�"�k���=jrv������Z��x���"C���J�C��D�]hB��o0_{�_`M�̲h}�ȏ��v���{ᕶ��X	~������iꄕ��2r�uW�E�V�h����d�e��]�\���
=�7�Wh��0������݆A^����LCd�e�i�礘W_�ɩx�LH��N{-�/���س�X�e<]b�oٍ��ܷ� h���:G��3u�������$��v�Y��� ����6jq!�"S)�x�qҏ��#�J�T�
��~
��AXz6 �#�_��qj���O�`���(��BuV���>�}�,�DqP���4�7z�����۩�&�w����)��YM��
�9q�՛�n�����H,	�	pT���'A]n��0R��)�"�bmj���kB�J>�ᱭ鿀(�������'��hj���*�c)��RHE�"u�5x��t��R>�)�q�< '�\`U^2��]��=�KA��+���7��A�Z��dP��P>�e���f�~�g׺CS�h�X��5;r�jD'$H�,z��6[��*�,^6%���:GsX,_��c���P��+W���
�p3R�w���f�H���g�+Am	2x~�� w��'b;]!��*]�k��fjb�V��Ǣ\MK��0%��E-1[���B]LZJw`f/��D�VgsA����E�\�7�"6H
C=ć(�]��lͳ��ZW)��6��o	,p�-^δ��H�+�b�t�?�D��
�7��u��Q�ZVo��t阱�SD�A�c �%&B�Bm�)-�	��ȢJ}�S�a��wh��ʳl��a��M��`,`_>��^��H���GO0'���_Q fKf6h�#zS�G��?�1 �$�ǈ�]m�7��ClR&H��r_��ʎ��DN4�_��TͶzQ�vh��/�q�q�05ù�'� `�ݮd��E�Ҫ���)W����>� oy-����9j�p���"�t\���A���u��V+�(S��������d��6�<e�b�RjC�+�'����[�MV@B���0�p݄�ۉ��[�1'�<��
У����I���嶇��e��R���4�M��=�0�(�Uݕx��n�n��\]�Gt�3�; ��d���?�<��_�~<�_;����M��8Idp��p��ڟ��ů����@��ow������J<���5D� ���m�&��{B��T��Ţ���������p��E�Ȃp=з��� ���v����MF��Ee���HH�C��2��Cl�(V��E��kaj�T�7�r,���RԠO��?,1x(q��x��찶ݱ���O֡+]�)��Z+B�����*�Юj<dU���Jc+Ϛ�w�K�P�*@:YOؿ�s���`N�8 �[�:�`i~ߧ�"%|���uN]���=��>��WZz0�
LV���5�$�Lv���~�w��D[�[@��+�ʳ�
lu�����4Җ .3U�C��	��������R ;���e��>�S4?�ܡ~�!��������A�G�/�>�����P�����I�ǜ�|�Yx��W��������eշ|��rÒ�R���	���j>BQB?����A_b�6 �dd��ӛ�r�b-H8����9�Ĉ�$�-T�5l����x��q)�=��
����?`1��J�Bן�\-&T������v�Rm�W�1�Ε=|2Z߭N���`�x�aխ�"��\�'X��Ľt`�~�����{�&���n^n��/�m<O�)Ӳ�-ua���8Ȱr%�_c��W1�Gis��)���H�E�[s	��qjA/�qLY��_�+ߓ&, 6o��U����(���~Hk�����`�!����N��nn���i�(���0$/qY�jb����AS�����v�N�~pl�+F��$D��ù5��!��ލS��u���*���75_T�+��*�ɀ��@�BP��?�(]��U<T7@��db�oR���D~��bo�Z�o`��j2�����mԢ?�Ag7r����^�o��	���m��͊�^sr�e��b������p��wi��a�x�]�R�0�5bIj�̆���б���?=����y����SK'ջ�$�'���!��T\�����X��)�ʁ-[g
Gը2�hC���O�����x��	�eۋ��芧�W��@�\�YV\�Z��K�wR�%�;���l	S��r=�y�J�q^�c�Q�V���M�f�5m�����@W�Ck�Yxӳ��z���U
���cn�{�.��~i���Q��G�u�t�}�=�c?�7�ؓ�WS4$���=�����owS�&�񞀘��)�j>��b(ui�[nx0����@�^ �]P�������u���@b�A�j���n���C�ɀ>��ݶ2FVϲ?����0v�yE�Tg���C��jj�����r��_�������+��koH[N���v{�����~�6J��]��w(�q$�l��D2;�O%r[��9��J|ڐh�ǈ����8�	�O8��Ȟt����z�8K���J�ޔ�6�����!�\�8��%d+c�dd� ������8{�)�^��lu�S�$�w92±�M��1q}ț��V���1ƪS�n��f�z!����ag�I���]-~��s�vQ�y�rq3�ᢘ�6q�P}.u��Cqj��=��f��'�
�|�9��mܡ�u�D^��:ߨ�4~z?l-䱹H�'�Z̹.��Ǹ=����3�a���Bg�"yp+�hbs��Ǣ �9+�{u�'ap�����:�@C}i+��N���s���Z�T�t��E��Wa
�o*�>~��GrA%��1�����@�D��Uh�1��m�z��x��+��o�Rku��E��4Oo!�.|^�Y!p��k�*��)�k���#v�*����\P}�|�g�5�'&��IN8�=/W3����"Pfz_�ơ��q�|�?o��b��i��9_i�6�2%w�#��YD�=�ܜ���sI��#)F�}���Mj{���ն��)T�5_@���S�����B�����~��G�+��W~U�1�-��c�RWu��K�l��`�o�*-MDt�*�F�e��Т]�B��S�Q������r8��=���?R4�Z,��ֈ��q9���C�yh����^�]u�T#�I�k���ĀP���㟢=%��ut3+tY����mJl�J%�L��;��k��%D�G��2��;JI��Z�,��y ���~	H�1���!�#�ō�)"c�f�%��0<����O��vW���gi����["�D�����;ȮI�Ʃ鿾K����I��_�^���f��Ⱥ~2Y�.�gu<E-)�i�C��e.�9���w����F��"^sJd�ۤ��C�W��$yf�Xܹ?��� 4#��b#��`u��]g�1S�;:j@w;-�]�Jl;oaB�4~	ʬ�	���/f���^�(��#��-�A���y������Ͻ��gE�[*,l[��Q�u����0�4�s����6c����a�����1��(�S%���v/�+@���9�����8�QW�Rv&pԱJn)a��pp;z2Re /�,9Td����{Նj�ɐ���W=}�b-,�l���-{�_Y5�����gt�uX=^Xo8r\7R6��s����g}����%͕��0%�"�7c"�Í6D�nC��8�4#43�v��_ds%OU ��C���~y$��K&q�~*Γr%��p���w#*+S Lы��uM!� :����L���v�}��Dx��0La�xnY��0%9Oa9��N/xߓ����A�eZ�����w���-DxZ���A��ov��"�L�\�!���9<�	(M�Uօ���sC�ݣ�y	%8�ct�u�ưjO�FTv����(�x�E�+�Ћ��|o��Z'���z㤃s��#.^:�*��Rb`��c��s>��3]���>���:{�%�j�.���0��T�ZZޢ�b�lEN��B�<��DA�?߿�o�*�P���N�@�'%���N�R��zWt\�S�_�{x�Y99����!1(�jj�1[:�
����� �B�W�NI��Fi����N[�W�*"�EAΈ�f������z��pg^��p3�����F�'D��{�����S�輫�fg>�r+ԁ�I{S�*D<  \�1�Y����ͩ7��2�Ll)������aPr���]��O���f����[<v$�!���.�m��B)��ϋ���x�CY�R�S��n�ý_�)��M�c��T�Tz`5e�{:�W[������"��?yG/;?Ыy�d��7*��d�`)�<f�t��-{խ���^���OS�0��L�3B�s-�49u1���N�x���H�
� AoU<���?R���JG���>I�h���@�����\�j��0��̅���[\�)����h�� [|+�Z���p� !7��Dw����*�}V���7#7I������kO"TB�藽$%�|C�y	 �¶t|��X�L2�@)+�b��1�Nt�h���7g�	�h9h�.�z���k=D������$�U��۩����4B������o�A�OS����DO�\ͳ���N��URl;Yh��}��Y4�8�prU��&޹F��kYmcbO�����:�8�S���Ia�j�uPnl7���	�{+���M��� NT#�J���FHQm4v2�����墝:;��>�- J��/�a*�+mvO�5��}&+���ςN���ԩ��*F�/S���,��:..�h������D*�蜒�K�9��ft���5�2���]�b�����b���0����Q�����$��w�EC�4|���nJ��˻R=����T3�L*�rM�3�Y��$X��zc��R���3�M�__:��&^����s�oC��}�9�R�d�%��Z(f0X��t]zۛ��j@�}X�z�@�i����7�D}%g�M/݈)��iU�Ύ[z����M�R�}�P¸��V\��i�?�a)RڴhI��}�wd��s@u辢ĸ��h�wV!s�&���?y��(�������L�I��É`��Tf&��!�C��WT��9��*�>9�&,'�$W�r���� ��1�f��q�C4C�^�H�{m��#��G���XU��D�����b��>�q��1q��3�zY�l/�7���e	�J�0�B����xF-z~���edAF�����n�T���h{a^���)���K�6����t�Y;a�>���9L�`�=\�]gN�pq�槙�	SR|?�e|ר��(wH`���</{��S5�^@�h��#m��[|M6L��TA$�/�_ ������_�RM1�Y��}J_�`G�G��@h��,�/C�U�)�(�*X��i9�v�UI�v�м��eګ><P��q�>vt�5�� ��rLm���,�	��em�iNBd���K�j�B��Q>V��*��|k�z ��`�WtzJe�����F�7��~_��d&���n��_��<�
wD;O��/��}���hw�
�g�Ŗ� ��1RhR� n�ON�IB�4���~
s5k:Ǹ�z�չ�0�.�Q���P(�;�+�:N@>��f�^QH.Zꈹ�i3K��aË���h퀂
°?�gf�n�Z�^�:���B+$.Nnb����x��9������%4X�AE��
U��bcό�r�B�f���Z�dF�!�pD-������v}�
?�!�����Q�y��a�w�o�䵍���D�Y8�jw��R�Gmg���k:R!if�Y���l����2�����Rϼݬʩ3bv �!�ل.5#Au��������R� ��o0�#�h ��x����K���z{呱�͙�?����
���0���
\hvp�~4{�٭}�O}c���~�jɜ��[|��W�-��[��q{�'S�iJ�8���	��֗0A8��{�����V�|�k�m� �(8��>dj	��AH��)�I�}�w��0�=���K�Uo�+�}L:*�~L�u�w�,�4�}!{1�!h��L� �\��kc�	���|���d�_8�-|lK�p��u�=9��� -6󞽒H!]OcB���J�*PgT��
6���VG݈�`LA#?��L�0Q�~UĀ����HlK"��������uv������e�v��	
��d������7l+�p�1)gݓ�'��GT��)2.iHTݥ�=^�\�TaS��#9׌��ѱK+@������wC� ��r��t����ET���?z�Ǘ 0%k����z 	��`��l�>�y"e���p�0���%q
јN���ɳ��W�ǲ� �����z��b>r� �ZЗ�H����n@��d�a���٤�O�k�`6�K|9�/E������9�ο�Ha8Ju��Thvv[�EՂ�V�/J@o��&G1J!q8o��:��(�� �`|�F�m fz�W�D���dfH:�����U�Q���4�f�Y��!fh4n��M>4�iZâe�f��c��96Y��A���;�{�Z�C:��w{]��ѓ3f�b�F|�G��I�q1!gOɈV�Ҵ�;{}�%�L�M|ZE��[gp	r���*o ����g�άfI흐�O�6S��r(]a�ҽ�
U��́3��,4�T�jq՚�)J;�Y{�lQ	�2$1$ܪ��(�����u�x���Z�����;�~���
[�sB��2#UR�
�m�*\'s�̂QH�$C�K�W��e�K@�  �c*�5}a�nv�l���ܨ��F��Am�Y��+y�/ˌIM��]�9���"o#�ѓ���R��rKc��j 
���>��q\u���B=�4�V�?�cZi'7��x�"΂����Pn���&n���n�R��i=��C���o|�]K��~}�Mi�v~�����c���!�9�ķ+�����d~�8�e���f�Q�,���D����e�G����3�1_��񻹨U�4η�9u;U�U�ٕ!�c6-��O��&��aD�#uf����#��!����(IPP���p��;�x�^������˫1m��+�T��w3���{A7n|�<gқ@��s��rc��3���ie���Z�����:m����^|Ͳ����N�ꬪ���"I��1	sG�p![�x��5�AoE����Q$�����[�%i�`�%�.A$�4�5��� �	�5�×�&�=>Mn�{&p��PZSMBhh�0*��+Û�󈋋Nf`Hi�;�'zN���D󓈥�3/[l|��TE�4�ۃ�'��%��J�/��[��jW?'rII��D���G�q&"ӏ�c[����Ӡu	�m�#7��z�fAZ
��h��
X�q�Z>g��,y�q�՘O�\��ûo�� vQ�CB1]2"����K�����,�Kj�s��E��1�MxA�6��������Zo)��t�p�5m�.��l�Q��̀���ī��aMq��bh���3A�P����T�=�]�RZ�>���h��� ߷�3E�_� ������+�F!͘������6B	T����Һ���|��>mz�E-v��5��FJ�3�Vm�T��J×L�I[.��+Uks����T�S*e�j�	%���2�у��G�1^��&Z���/N`q��G�k��cc���1ԙ��a�/�-T�h�nR���W�`1���馩5�1o*��Ep���b1������t_�����	H���:�����+��˾bD����n�7�K%4�w�η����O�a�5�.�e\R�D~
��nAI���y��� ��R�b��eȸO�\��M8���X�T�K^�����������T�g!�O$ˠ31RxG}�)B3/�d�2����|w`���7敦f=��͘�Hp��2�8�߬�=d���#�V98E����� |��M�P���X]�PJ�2ꤱi4��҉l����'^.I���l�^�]>ǣ��'�T{��h��V�@�ֺ�6�)jq�ܹ� A @��������f����1�]-�1H�aY���i�.M����Q �C9���Դ�"n�Δ<\��0nU�*Հ[Y2�}���=�k{T�2�`��+c��t(��3,]�~>PE�#]Q�B̓x�X����7�/�0�Y,n��g��_u`�f�z����VU����t	&�c+��U6/���nP�]j���b/E� �:�5b8�5%�!0$��RWPhx���Q8W��&�+@F,�`�6�ĳh�(�
��� ����+_˹�;t�W-�p;`j_�>�~���j�1¤�,l}�~%���L�s[�aX�)��ja�FQ;��eJD��+���\&G����r�bDw�z-0m�2��˳{k���(����/&'-7��%�4��l0���)��(�
���~���c 5P��4�*_g叼"�[�,�VR���L�V�%�R������<7��f0q����Wd�:L{4\4��XQ�1O�9^�v��f��gQr^�=W��ދ�c�p�J��QlPC9k IhD�8����3K�(ޓ�aL�N*���+����2���g_��dg�H�@G"�����0'T�)�֏�23�J+�6>����n��^����U� +i?45�² U�9ׇ��8��������]@�D�~�D�k)�\�=G�C�Z$�p��25���E@>+�����Q�A�~<���n��>��l�H��i�<��q�s~ J `�'6}�\w���m���?29�	 
F��3�=2��)�0�^��c{~�����^�;X� �o���|�q�&�Z~��?��:I(E;�n��~��ͦ�y*��3x�_�P�
[�\�4Y��^Ba���Y�EzR����]��L�da2)o���_/��
��5|�����9�!�7>S�`���M�Gtn��ﴁ���4ׂݚe,RD��È+�XS��=�j����a)��d�1�����mT�!�5O%�'��\�����������{�B=��K`�I�M��&�&�Z��O@��!���|��O��`p7�3-�(��P`g?����p�S`�ah�L龻+��qc7l�<�����`(���M��.4��Q���y��W_s�}z���G��J��ؑsu{����θ����B�݇<�Q{��2R�I�fg2`�-F\H'�#}�Sb�P��B���6�)�\-�����2[�~hg=��8�I\��i]��/����s�=�ml�]��tY�_�����j�w�<g���؄��:|\�?K�Y@���>��6Q�-�%�z���݈�����+ �3s��N���+�O��ܬ�nZ���p���r*���\�:qM��:-ܬ���9O�)>�����T� _P0����n�gW$�Х�8j3��P��C������W��W9��p�:�b�J����)ד@�T.8���>�@\��70�����d������XFAB(���H��P�
/�C��KͥU-SUt~� D~�U]� p���%�)R�vn��p�� ��(���~'�]���B�����q7�W�����U{a���"���aGCX��*�n����fc��4���QWI;�d2�����ݚM�!�M'Ǡ�$ƃS��!�#��r��Nns-/%(� Y�!�l�'��+߅�����v��7��WS��U�#��o�>3L2�CJ����g�Å<	�Q�K��P)r�Č�I��t��'z�B1�m>w���Q�VV�뒢� #̣�l��������-�J�L-�e�WU�%k�d<��n1�j��$=lvB�6܈�Qbŀ&���\V��VM��3 �[m�Ƥ���;�e3����
��-4�=��ç����g�$�1���X�u<�����Z��}��1J�\5ꃖ�0��������k'��$�`���O�ϰ�K{G7�|ࡓ����m�i�T�*J`F��W���n3�M�z`�di���}�3yl{��#t֪WX�}�SO&�3gz+�w�
Iқ����,����DZЇ����ܽ}�*µ��[�݇d��D\�qr�1�
���mKz���9[Sb�EK���`�^�z�5W�〗����ν�(��#D���SV�nc<�8^����œ)rW���A#��W)5 ��m�S�:�"���. �1�o�c�◺��+]���K��h��lr�{7&�-�AU��|8h,������;�S}����oB���F��>X���N腸f�����C%�r��M1"�(�_��GM�xe��(��`�@�����v[��}�q3hC���U��PG9�s�%������ގ��(d�h�PPM�dTMR~`1f�m�
�z"ב
9��� �I��z�����SG�.ʪ�DQkb���M��X���eT>i�qf���.��rJ���LLd�<� �iA���(59�����Uѕ�eX|m���/��<���D6d��^-:3��S�
9TJ������{�_n{R�7ѻM��o����������ѲKT��+�O�3�Wŏ���V�3��t������Ϝ5������:k.Y�Q�!�WPX�e�%�ƱV�G��b�-7�u�H��؄�x��ד`
�ҿA�ߦJ#�!��?N�֗��Չ@tr�e]�����J�g{'bE�<��� 7s*y�<e]��%��V���,*�|C�����&,�M�t�7Yg~	Hz=�~Bv�帨�Js]��m�h�vȯ�g>�6%�W��;���5��x���b�T�y�������h���hw#J��ʧ@y��&,��Kl�Y�.�P�_�(��}C���\�S\g��~%�IQ�����+]_�&����w֏�� ���2v�T� �7������J�b`~���9��N�)�8���Q����X�+��m��5%S��V[U$�ߟ��R��Ƕ��&e[6�L��w���`�=��O�]��u3I^(��d���|�9S�.�P�gx�p1j6$Ć:3Q���� ���J��#$�h ��I7}�9u#�����3f$��I�
���ߟ1��(ٹ����X��9"�)Pr��In�/�o���X���J.Zp�bu�R���^�	%VU=C�3f�����VxG��ϴ��,��b�?q�i�/���w�NG�Ra��l��~�5'�§�O�����r��I�*��#���6|�no��u���"�;+���W�b��ׄ�t��i�>��~���/puĊÊ:�t�;��6?������ v�
ט��<�]k�eh�8�>��� �.�gA�G�K�\�%R����)�e��$�j_��{hLެ�j�������U�]����C��o���c���K^��-g�\��$.�d@��V2s��J�ړ�͈JI���|��
%i��Ǩv~83��N¿��E<5L6���u7�iG�o���� �s�8�|��7[�����h���$)s\>X�˰�~�9�i�&X�Qs����𧎲�KI6a.�����s&n�_=��QH�'�{���6j���z/�k��P�k���q��4��'Ri����7:��h�%�ҳ���	��_�FP�ūc�#6�*�\ځ�*�ƯYQ��YW�CQ7� F�lM�z����w�8�Eo���Ğ�8��pŪ$����#H�q�0N�+cS�����;�`fm��rR��_��,�q�BX��w�
�Ll"�|����]�q
��.-_�-ΗV�[���^������6'.��(�L�N�i{*t��S��p4�	\�3�6ξ�&�F�����4Sv<��u����d��w���[�h�`�[P�$RP�e�Yf|��c����G��4DG�h=-����7��kU>��0
���K��g<�kB��ީQ��$�lf�Oo��_K��}z	e�������9�"P�gFtT0�FI�!衢=��Q4�����k`5
�B\b%yHX�#D��T��w"T>�����к�Nyυ����My��u-HB1�:[w����h����P��o��>���0�P����Z�Od����5��!�e�к��z��[GA����Q��c�\�\�y����_��2'ɏ����Uu
qg/5~rSYqxV�gZ]����N!�}�p�ADm�%Sd�4�)��=����SX���]}B��B ;�y%R�11!t	8�V�=�����C?��(|��C��'��37���VB�+���~��-�I�ۍSCߞ�i����,�^]u�b�����@_�b�CQ�~8��+�!>�vuK>���O���<9����5\	N�[ei����?�/;��RɃ(by��A�8^Y8�+��M�����P	����n]g~!(�y[�^��0)] fl5�mHAW-�U��ƍ�!7�����@*N�Q��j:+��C�� �A�`�������̭����0m�_j���*D�!>D 8�g�q[3]�5�@o���`/���B���,�Z�}��G�z�^��Y{u\�/CBE\U���ښKϲU1}Qw�>���GCuH2Y���!o���XƗ�Y�Β��r5yq�d)�(Y�������C�nn~���S%`��=�*����U�C��O��;�7I��H��G_����p�[��8�N��4d�OF�E/W�0�V�.:�<��[�o兞� L �����GZ��*�:gb�V0��K�<�qT�\YŝW|��G��vx��~�o�'"�_{�d��Z?��e��f���U���Qf�s4���;�p�˵ 3N�b	S�5$g�
�;�����rFB�4�	I8A�@�B�i� ���6�o�)��k7��ّ^WLk��;o�I�#���s��Q�������N:k��.5-])��7�'�٣��r����c�8��*oWtL�2`!��+]u��~~�.e��Ua�AT����cu�)�nH��7@�"��ݫ��y�gieM�	��L<��[ʱٸ������x�m�W��Эqf���_�����ڜ���M�����/�ؐz�y�*�<+�G�����O�����)�Ք��I�q����Mg���O��k	���PÎ�za�x�T���"�'�%��GK�g���hp�o-��dHu��������A>k�g�h�zm����N.�ء�]�����NA�87�bE|z:�]K���C��Ğ3��#w�2�<��9��,)���xy���]Lnn�A�ͷ�,\��Մ�t��p��
H��-��,�����LﭱaFg&��?�a�3��C��������A�)?���A�<�$-K���.��(�Պ�	�4���d B:��ci��}r��A��C�&G����te��@�,�[RO��5�h>C<N� �?�j�RGA��?�^mz��᣼�t��{<�9�Ơ٨�9����#�A����9v��a�5a���MF�+��ڙ���&3�;'V}�/d/���H�(�%P�X]����:S~�g��;�m�p[���(��˛ݥ�k��B��6��I�dZ�\h�ĴJ	������z���P�|I`��`��;a�j�*�鼂Z��?}��|uV���/+6�qJִ���x��������Pܟ :B+���)ȨJ?���.^��� ���S�o���7_����/s,�}�p���1�4T�a���Mm�����w��"���������:Q�I�sk�i*ǽ; ��g��fyJ����� �Mt"�/Y�=	���M9 ǆ{Ϋ����_A~X�{Έ����������ߓ�'C0��N��9�n*]=�&��"��U�m�[�ܑ���Ԕ�w$D���O�Ԡ��\Y�w,>]>���������*P!@�C�7{������'t�c�D
�����B>Y+��i��aG���� mtf�(��q�X��?m���d�m��C�w��d|UX/L��I������dg\��}v�Q�1��w-�~T��l:���8�/�=��Z	�Ҽ^m#=#�t�K,���6�]�q2��@�b:�s>�<4;>�	A��p2�y��Ij�@�Z���`����A�/�O@ �ƴ����}�_Y �h��R#F� ���W��0K�f-Xt�+��"!ɼ�lV�ͅ���Z3V��}�P/"Oe�J�h�a䦏��8�^���g�������߬�#7%������~�KW:���7�u_�<ȱS��SPI`�2���[�2�Y������,��+O��ʡ��,�Fߥ0Y@X��AC�YA����g|s59sdHļ.��ר�Ys���9��9��[�Y�ӅU[��E�>/�0��-�����4�xF�P#J'��ү�E����Lq�2����mUI�� 6T{�Z#�����3Q��Q�砒�nj]UP��$�����A�޻f�L5�钠V0�vft�@@�v~%�@
�5-m����2��?4�[���	GA!�F�lރ�Xc�{���������Р�Į�혷P�a��v4�Xco7���[����9��s�$�_� h���TW�(%�G�=�&p�CuAAr��;`<���� uŹ��x��y���2�r�
�ɕ,)#D��!R:� ��eG��-S�{��is'�n�Z�|�9��Mہ-���ӓ0U'���_&��}�6�Ԑl��;��'�J:�8�P)�L��U�a���@�G,X��Q���x� �{���V��2�<� T���ق��mح�:���Ru#豒s��Q�=;���*6�U&�!�{�-Y1)����b"���ǯ��+�ė4� P�r�I�.�෵�5J�����j5`�H�h�(/�l�`��`祬�f{��z��?[�^�Iϓ:��0���0�K�w2���L$�#�n�nw�P�H'��q�m����$ԕ���בI����_�5�6-���8e��{1	�x���h,o���4����K�t��Hף��t�Fŋ��$=������9��S �;&<�Ic�BV�0� ,���X�{���>��[�s���-'+���0�b���OI�D˧)2�����*�OŹ�2.g�xdBy�q��ju���p3��;a� �.;G�s߭��;���f�X�i��	y��KI[����z��I{`�VE�t,�<�zC���ET��.���PьsVO�L�~��Y�-R|�7@�j�h�oG��_k.��MUw�{JM��;:���4ձ �i��
͚|��刑ۮ�*է����f\
�HG/�Zy���FQE��FG~5����
L����@�jG�F.�U]���UM/�nm�?��S�W1Q�E�,��>���4����5? ��7���j��I���4��78��.z���V�y�s�*MP]��-��[��-�
�����6�WHS���9��0�b�Y<n[uJu��M	��~@	����=�ɘ�1S�Y�"q�\��`$��`�6������[��?����d['2���|Z�  .Z^�k�L\I~��`���*oq�8�Ċ�|��1.�=�C�^�հ{�`�/�&,�ĊcQxT	M��d�.�/Պ$��i�F���&ӕ��\l{�� �\>�{�"h����oh�k �iJѰ�颺�iz՞��B�OD �c88�Z�w.k�g�4�7ۗVj�#/���!Hn����{,C�C��icn�|	�9p�S�W�������(zb�h�T��b	�~>ߗ9�z�P�;���⎁�:��rj�hF5�3�&���?��yK��!A�3���/���"o�[Y�8^���>)�;�MM�B�&���B�6jk)$�4j��G����,�:#G���;� A����������(�Q]����|ǳx&W��e���6�z/j������
$6)�ѻ��JL\I2��?��o&�%RV�i>e.��3�Dl�����\�0�0�!��m�C�ԣAq{f��\,���L�KA^������	��л�ۃ~E���bIPYh�R�.�I�4���x��66鳚ڪ�T��j�dnQ��Ж 	�*�"Ns�m�Μ6/8��$ds�ފD��P�+������ǰ+h��|/.��jv��;2�k�߬LT�̔5W��j�>��'j/��.�FO�p4�*��;�n{ A��_�oV�pL�Iy���e)���[����%V�p):���q��$�J��"��/BA����I������`��j�D:�w��,
�pGY"�R2����ʶ�)[���zG�2�WYM���klr,�^>S��s���>( l��	r���4�ٲ�>�:����ϱw8L�;��� ��|uX������(����#荟�0��r��Iw�l{�2�M��{@܁�xH֨c竷^�pCY���~��n�[k�32*��� fe����j	3����|��)�|H����{�[�Wh����x�C�bU���)�;N�E[�'�;�e?ڍ#Z�K��sޖ�4b�;�Y�Jt���[ԓOl�EG��H�l��gg�8y�U����~{߽���>�_��_�'�!��9�M M�����p3��S>����51��TÏި)>��i���[�^:rA>���h�B()f�����<�J��1�$��g��'�Ϛ�"gkL���~�V��P�~u����:t�#���{�����i7/�CҘ(���M�U@�
l����Z��`%�6����X;C�@���M���p�X��^�ؑ�<^>���ph�eTaΥDo��b�]]�d�9���VB��T���w�ѽh�[��N��2�8�h��]o��W���>��%|���kL��Hዠ,�����j*2$B�Mh�F==o��ʱ��m\Y��R����i"����g�׍�CG��`�������fi,8�}�s�����5�7�z�6�w�..�X�".e11�[{ks?�$̺{=E��\�e_���(����S��K�o\�yNHډJ���:�a��1�Sg����/�ѕ�I,�@�x�Y(�W�>?��SOk�C9���w8�2�6�n��>&�7�[ۥ�X��o�E}0%�,`�Y'1�`3�ٮqҕ䎦��2���(:�
=�0�Է!r>��M��[�v�^�{������&{L.ϏG��?�)����	C֑�z�K������:��C�w�9&�&]H$�W*��a�6R������&��8��B�1��}S��C��+)�ٗOI������O�4�k�� �k2�6?��34:�r�V>v�k�?�D��Y�|�S�e�>&9 ��z�WA:��]��`��@�C��Q�AS"��k$�T|<Apo���\j����	���uw0l��槕�C�9(�u�Tm9��w�^�w/���e�#����h� I5��r���O֡�9J�(U~�c��s���9�'��ˤ��K�ˎU��y��-n�C�D������J��W2���ɒ|�`'�d�?ә�������*�V�����Up019;�Z�q�4�"�z?�4gz��EY�uY��βE�4U�[����~��h�{��2E:�`����9����F6cl����,o�[��������\������	d��"*�����%(P�o�0[cf���%�*�@<s$;�pb"uwL��_�-�Qm׽�5���(��AI,6H������	__�K%�]��` ��3�V@ �:��s&]�'�T=t5롔b7T2N��`c�Awv����<�3l�ZJ��f���%�}R�y�� �h��d��(��l�/�&DwdL��C�NK�M�1�KSf֌{��fL������1BSS�X�~>�}4�hJ�0�3����B	�ؠ�~6��j}!Y&�P��:�`l�� ���\=��)���4�����zCb���'����Ej���GE?�K4�A�����#c���ת^F��,�dv���?N�CQ�4�Q���k2�xCRzoGE,;�ūC�3 ��`|��h�~��9�ů6��R���*͵�r��ڒ/�d�vXqC ����w�xuq�)�<��J�k�:�(�!��S�����:_�Y�-�}h�����N��ӳ���/PH�=sG�_TL_y�I����-\f�.�g���n�"vw#�g��L��kHИ�5F���ДN B�XM'���C-ʇ?g���M�n��Ĺc��7�m�B�={d�'������1��p���J�]����+�`Z_z���	=�M� ��+V�AˢT9l�)�d
��=-��AEV6����͞&���}	Y������� �q���%?�YR�~�@3̕Ys��-XA�&�윟XǗ��ٵ[WŊ��X���&��F0���iq�
S�Y*��8T�����(��>�-�-�>:T[���76:�y��c:J�<j�Or!��lw��	:Ro4u�z��I�	a�t� ���ޛG92��l�c��U���T�:A���.1&�JM�?�*���D1��C��ѥ e:��"p05s)�Ϊ�5������#�椐�6��<1���&~�S����ꙡ�	��:��d�
9y��j�F!?f��[��tJ�#W�K�GT�'��(�'��/�}��M��.w��;����x*:`ܲ2ҮĚ�}3�XAR��l=�@��Y�~��I��7�C^��>>����FKv������ ��6� g�)�[9z��"ï�H�\���~�3�'�j_�,��Ɨ���c@��n�ͫ*��AEIT�u0,�!��K�!��>!�sK�~?����RSK*|�e8z�qom�yb���s(�]�-��-��vE_Jd�q:��eJ[�ګ�`q�v1�@���Cݛ���{\L��~!�9��ﻧv�)���^3�u0}'A�N��Ճ>%��8����2��"�o	�xO���`{PAc8�I@�{�&f��)GW�&����!QзHc���9�.!,�����r������1	j����M%n)qC�/���
 Ua��u�*hLk���Z0?<�a���W��R�%���w!s���0�靕���te�ځD�z ��X��Y)̇'WX��n�Ѧ��>b@��%=����z�]�U���/���r���ʽZ�k�|>�+wӷ.�x��v�n�5�
�I���V^���m(Z���_�Ǘ7�d�X���Z:�s�.�`���9}f�)M�f�K�Ιe��mWވL��Y�ef5�~�T��ͨh#������ujz�*�9Q{VȲ@?�+�Y�al��}X���#L��H�1(��U�p�!N�ۃ&Tiw9�+��Hd����ќ�����9W� �G[�2��(�����Һ��۔� �F���T�ɆC�05�ft�Z4�Q���x}ղ%K+��S���#��<��9��.�['�D]]>��0v�=��&*��'�>�(��oH��O�#8�@#�Uł=�m�g��Rq���8mum�D���>�i�tw�_1�l�E�.��j����3`����l�vջ ;r����֑�#�TJ�蔮�n@�<:;'2ߩaZ���rb��J#f�C|�7����(eD�}�����E��1���UoLx�7�}*�����$u�B�p�.X#Y�׿v������x1��w�?�=�H����B�Vs����=��0��M�r��}7%ȡ����9�,Qy�"���H)��c���<��� �Fue
����� �e���ÿa�^;�
�w>�������t'@�G�u��hQ���y�b0H�!#�i�h*�c�u��$`O���RL�a�C@rr���ςT��PMQ��M��K��+��:�#�ZXnrz!�j�Z�c@zp�؍�[>�����|��m��=ǘ�����tN�P�_���W�	����oX�(T�.�e�$���E�?6�I@$��/�д8��G~�C"x]�Pi� �L��� �Z:�3MF�����l�KJ}�|'�QrY`�X?6i 0�"U#��5M�r���
�1r~"��2��0�[�������D����5�*�%=C�1U��q�˅�����w�ן�o�˗܊ԭ�	�*�3���c����,�I�����]���W1�\���d��S��i1P�`o#E�8\��.�%շ�Yf?*�`��*�<E� ��Y6�g7���kk�CF��"� )fK(�g�0��ݍ���U�\��cH̜���M곝Ϙ[Z|c+���D�n na׹nF���HQ�l�7^((*����Q^�i~\�:m����4c����96�}�q��������k#�Du��>Z�h�)��(���������M��Xx�g�Rꉃ�$�ZB�ίzj֩B����[U�
^p0Jx�@l�!6�.:��Uނ�9"pC���?^�5A����Tvf��0}��U� 9��Q��8 ���^u��52� �jͮtH���G_ym�0���(��"���}\e� ��X��yI��>���O�x5B�H�S�
�����.\�>��9��ٿ��g?�7�ڃ`��֪��C�\�qwa��{z�C�MP�]�\�j��:�I+���� MeR��f���,e�=��"�f�w�ciG����j���n�9L�T�q�(DP�S�&7I8�EI���`5Eb��Y,�7�;&�Y���A�ê��9<I�Ͷ	����!��Du��^?�����hm�܅b9�Yzaq���À$t��cȾ�N-='�/����EU������.J� ٱ��%�W,^�7��h�����я�e��La�N�bX�*_"$}(�1o�=p��=]m�Pl�P�$xCt.9P��w{V�7�2{��#��t$���o��l/�8���k��&�5��Q�Ͻ�ϬL�-��ؤ���rƗܑ����h����E���e	P���lԀ��9���DI[�[^x$�o����eŞ�-���ۧ��_/1c�Su�g�ړ�B�j�Yo8c2��z�omb�&��ӫ���m$���2�lT�,�{v>(��@2�.�ew�T�:d��j�d�1���$m'�p�EY���Sa"S�^���Y�ɴ9�8�ig���Hj$�;-�+��l����Io�1p6�0��k��]v���$R����fd�O�.�«�9�����k�2���y��0��{]�8��F�W�l좤�u�po�L�=���i�"y��_��&�1�I(�j� �����[�C3=Z���,E^r�R0\���$�:�j���C+��������,ߟ_v`̋J�="ٸ��g;��X9�_#Rϭ/]Xi��� �!\�w���z�v���:�̪/��4����Iv��) =�����|�������!Re�f��}�b}#n|=qb��p�x�A" �E��g���.���S�珃��e�dA�r��ě�]��++��.@Ub��2Z�
)jER��貭B�cG�����D<C��iF�u��!NF� 'n�G��%L�\SP�UA)���(�Y=Ӛ�&ZH�+��C�4d�F2|Gރ�;�+Ӎ����͔>,[�\y��D��+:%�gL)ˊ3) �,�Q���W�z�$Q&�߻L�Ӄ('���~}����}bp8K��a�P��˶�!*���3F#���!��ڨ%-��3K�ˍr4�W�\OIa �0b��z�1����=
�Q�jhW��޲��Dq�)|�W�~�IU��r;̨Z��av�kS<�C	C��8�s�-� �P��5��Hk�L��6�BR%Q���
NG����e���MGm+�c��bL'�ҽ������xѸ��k���<puJr���-7���r5I���H�X�L`B�r[�R�5��jl�qМ�%ķ9��WF&��WE�̈t%��W�����`�2���⮝���M���X���4��Ec_M�o�z$u�D�%��-��?U�^���<����$��=Y���~"X����)��I�wS��V?T���C+�����rFr���$F��nL�	��i��C'�O��>�����yp}4j������@'����� .p�6��U+�׿�,�(1�k�>N����5�V§3����4\@Ђ�~)�{����-�2^�lb��?[�X2�Ig�w3&�0��z���LQ
�L0��nyp'��;~�yV�
��Z��P�S�h�-2��I�$K�%�����_��QL49B��D>�l;����=�����d6)iXXw�<\�s��W��0S8f7�F�b�ǧU�n���B���,����c����K�[�z~^<Z����Y��?��2;]���i��T���6v��î6sC�Z�mN��N��^l�w�%��}�B�5��W:�Q�}��Ε0mMw�C�я�דg�poj�,�4�AB'���� %T���?���UX�Rt�+s�s"�>Z"R����L%��@��Ω����{�Ι�$F�����(.pTJ��2�Iy���5�B����E�u~:lq1Ž�Ĉ��.$�w�vw���Ȥ���Sr����"�]Li�&U�;p�� ��l�)[c��*6�&MH����4��bA/��O�e_|Jd){5�a�Y���_ݪ��0%SBp�~�V��w����?W6��eT�v���ን��\�1���90[L��%qz���\�����e>�Ϥ|-E����FO˸yY��Yf���n�/\�p�v_ыRU�8&H
�t�D騢U�o:بU�(+h%ιz��n�����0o���՛k�(h<���㇡� �(u�W��少��)��P���R��f��[-��c�^i�޼H���6��J��{���>O N���q�(��.Y� +)Q�c� T�p>AQ��`����{��xʝ�Q���(�	�4o�:�gG�\�+`ע����J/}A%�n�Զ��5L���L���o 㲦ln� wfnp�k�$7���U�zGN�G�D���2X�n�'��(����ɋ�o�5�g #JT�Dp�t���}�H?熄�?��ҭZp9Ä�&�L�#�d����g�ݣ��,K�^Ũ-(�FEbx������A�-X2T��I�r��:�z%���D �ʳuz�9FT��fzƧb� ��/�"���" O��[5��Rp@P/�B?�T�	v�贄�״�b��E7B��T/w{]?��v^n|+���j���5��/���|G��a�t,��8S�.��I��΢w�hZ����,��χ@oA�<Z~���j�iw*�8�l��]�}j$���>��#�}Nr�=�����j�P��PN��7�b8��ݥ}{.��ė�.����	H8����r�M�3�.[�b�v���(��&�N;������ֲ��G�z��m+���<?l��a�3�1�)����.���ⴻ�y.�;olx�F�Ed�W���l��7������ݙ�q�c����-�8��'y"�� �L�<H}����Ӣ	>�c25\\��-�^�:�^���f�1�/�Qg %�x񿎓q������Nm��x��R_������f$b8%C�[3У"��rS�t�Y<�O1���u�q�$4�"����K��+Ĭ8U׉i��Gn�ї�gn@fi�p��}jS�6~T3�Ta�S��<{%n��(u�D���q�����`�	�I��=��o�u���O���ys�<r��Q�=P�]�]�>�*/;�5�Dmu�����;1�<��4��֮a1I���`"�4V�ccC~wT�����_n>S�!4��� �r_�8��u���\��eܒ��п�ax������v{] @m[Ibߡna�b��тe)������K�g)��۱���)�R�6�5�ʰ�������^��~�'ǒ�N�mE��Vz*�s�ܼ�z�R3�7�{�A�MD�`�5�Ĥ?TS���M�zQ�0��9���<�5�S��v�f��b���m��x���?9"x|F��>�Шg?pg#�H�X�R�����8����s# �@���H���w��8$��������Cf +H�Zc	���<�;� ����Ip�e���&������!����f�ex���f��LM�u���H�+מ�\��KE��� ���L� 5a�w�A ]�+H�D�ΐ�m��ugu�ds�y�]�~:�n�����b�	jt�4����Ƚ�P_��>����8l�u���۶!G!���u�tp���h3yA u�Dr��޿�'�ۭ��ކ��*�p����W����å� �yi�I����u� Ϸ�a�!^���5�=�u��b#�p�����ፑ�t�i�*de��|���~!R1�˂Z��jQ#a��P�T���4�ڢ��A���t|�i�[D���0&?���tȜH��b�q��~�t��|Bl���Κ\j�S�[�[�6+4����|���y�E�0�E?�Pq,� �C�gR�z�ro����HV�����3�%L�.�����Cq{��������1r�m�� ��C�=�Ƴ��)��Q��WQ[X��x�n�X<XԆ�[-���}��
�W�؁����Qߕr<H�_V���E�@�?R�PT����X�u�i1'y�z��.EVb �ڃT��SM���1tG��5���(u$�O;a�%�B�}h��(��`�����ֲ�|[g��'�9��Ԝ����U��RW��/�|yY}��#<�}�9�ލ8�_�[�eJBQ�?�,��E�+���6����B+Y����;�Y�HɭC��|�+���/��RN	1��J�Oi�T��~=��@4D����_�?�s�y��U��<�yI`�L#����t��y�.]�`ݪ���f��K�
!mB�j.�ɼ�H{�m���Ђ��^QfO~����W�@H�����(iH��D�Mx�Y�N�������t@'�ίu���E[�]�D��* qp���kRW�}��byꑛ��s��0W7{n��豥z/�]r٥�Lc���Ȋ"'��\���ވe!�T_q�#	i)�B1Eynٔ�oD��7������T*�pX�I�Ur|�Ar�lɣ&:���F&�;�q���΄�L0ǁ�����_�|.c~�d���ϣ[�f�,�1[��Ϊt���;���Ux�ۼs�Xv��P{��'V�Q��pȟ��z7+���ʇi��L��-�6���ey;���ݫ�?�썟�ʙ���+�6^'�kt&E��$�5�y"Ր��,��|8G�mۿ%�`�����9��h:(�,?"6y����ǅ�a�����Z��ʝ(�8,�9�̻�@�܋�<������� 6��慷0��Xε�V�=�j��.in�������`�E�>�z��]L�\��(�v�-CPE��k�L3���,w������~z�N#f.eD�Ж"����-�Ep0w<���U�A:?&&�tI]���Þ���y;p���Ño�l�:D�K����Pi��,5�"�~]�����������+]��y
1��XIݰ)�YN��n��\3��¸`��g69�n�1ʻ��Ha
i<0�e�{��=h���.;�Dpi�T�&#�3Ji�a��"5���l'�K�(��,��8ʙퟛ�?���bĂ�z��t�����{��*���� D���:�eȒA0�����T����6�Yh�I ��A6�<���g_�
�(V�5gN�bV#ĳo���$�z��=�f����ټN@�".L��D־*i��^��0�iܚ8������+�	@�=d2!��v�����E��W�G�����]}Ug��Թ^[�-�s5R	�O��[���[�|w3�R������V���[x��"47A��b!R� ���gG�EC=�9��u����5٠~�d`�w�쒇��$�"��p����1u�u�f�yLZ�~�s�ou(,8�U��I���M+��~�F��1��ɷ$)�M�9�Z��Q�[�JD-��y;�P�o z���xb�1Pg�Ga#K(��%W�̮�ؚ|�_˾I��/$���aQ^�оb9����B��Tv�9��C8t콵)z�ĸ_�F�	���6%��}�<��3�#�h�]��MҼF{�e �S��[���YͩC�"'�9FZ)9�˶��.��9��͞�b_�k�y�MI�0.�IA�t�=T5h�өª ��;���q�'��)���Z�$��,���8�J::������^���9�Z�-���FU�1�_t��A�1�{^i����QQF_Ks� ��hY�:��N[���5&0��)��J#d�蕄q%��GÜ6a�B$tk��*4��)L�fY�N榴&�kJ�x�׫�,\���y�Si�i���i ��^���
��ai���?^���ʒMȕ3���e��>��G���{���$x���|�*��0z$$Z���'c�m��q�S�rܙ*>P��~�!P-�De~n#�;�F+�5�M��[�����uj�P��k�
G�5:��,\*��-��,p���p���O��
m)�p	�zN2�
)íU�|g��#X�9,��-X��0"��1�[�\��ל��B������e_���ώ��(+fq��=����^��0�:9��lU"�_�Χ�Etx��[]��F�k��`�Ç�o��t���'-
�fa�6N�׸�_��lv#��Q?�����O����PJ��w�e'c,��#�߯K+���u��F���1�nB�&�Q�2��k���J�L����ݎYY��!�#�O�����	N��'SL,>
C	b�9o�e2p/h�+�"�OS$�.S�q�O^^˩98|���~����Ϋ>���w*��x/���:B����ԯ�F��9>Dـ*NR��k[��q:L�<"2(���^�,}W�'	�XVQWtZj��^�Ȗ~8���C✚�Q� N����$���K*::y:�����V�3�ɬ�	�����u|� rN�ߩ�L�~�&�	�������H_��x�d�U�Ɣ����m3d
��y)�,�k�>߹�:� �d��h~j�I����)TV6�^�D���m�N����j�ȋ"rɯ��8Q��Nf(�.,�9p��-�Ѯ�v9<�c狍q�?������8ů��|Ph?�r`�N�Ք�ܔ��Z#xbK��*]a,*�i�����>�u6���]v�LvP7�c��(pJ��Y�O��Lwm<�v�W�b~k��q�'��y=�?Q\�e#�g�[!=豵�z�y�\(���$�N����Q�6�_D��<���%��}��6��&��&WM�����)鈣rmv4���1���ş��V�#�돑TŻ����������J �F�Lm�i����zQ9M�M�2� 鄨��(��݃���<������L��bAv��M1��cw$릛a�&.�)��)�����F	������X�a��˻{����,CL�78[�`"gŴ�3�0+hB����**_��[�M7�O��́�9U&8԰G^\ Ԭ<�JI�t�#�&�8/��t�Cm\_>=���,�C��?En�!sp�B�d���g=+SBW���nW� @>L\�kCBO�N��{�sD����&����lV��|�~IIw�mh���Du�:W��>jP6{��({Z�X5���U}0���8�J|�Z��(��pɱ������Y��VZ	{��e�l�&�=%ty�̈�RP&�?�R��E���C��ƨ[_P�ؗ\Wk'Qĥ�9���ցN��	ڐqr��X|���v{�\$�?#DtxukG� C����hU�{:B��l㤞ySm �Eg�#yt�	�\)�S�A�9��S�g�C�|C�jLv:M���ʶiEh,�#R|����e���d޷F
[-�l�*(e8U�88��vM���?�g� �t�
;q*��:�4K��/_���W����n�m���a�׷����J�Y��ф)�.�w���6��R:w��m��1���Z�"J"}�?���,^ѻ~X�C3��Լ�nXX(rяs������Hط���m��u�%�K��3W!�J�æ��4�l��Y�qM��_�֩i���x���1��D��T�Y�~��z{*~�9>�QF���۔�5ET��{�R��n�Xؖ:|苭�ߏї?����{�)㞂T
*��8=�����V��n"����/BYUk�neh��e���l�wm׎_��>�f/D5�������>Μ}�ܪU���Q|�^�d%	dDh